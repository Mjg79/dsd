module jh_round_b (
	input [255:0] in, 
	output [255:0] out
);

	wire [3:0] sbox [0:15];
	assign sbox[0] = 4'h9;
	assign sbox[1] = 4'h0;
	assign sbox[2] = 4'h4;
	assign sbox[3] = 4'hb;
	assign sbox[4] = 4'hd;
	assign sbox[5] = 4'hc;
	assign sbox[6] = 4'h3;
	assign sbox[7] = 4'hf;
	assign sbox[8] = 4'h1;
	assign sbox[9] = 4'ha;
	assign sbox[10] = 4'h2;
	assign sbox[11] = 4'h6;
	assign sbox[12] = 4'h7;
	assign sbox[13] = 4'h5;
	assign sbox[14] = 4'h8;
	assign sbox[15] = 4'he;
	
	wire [255:0] L1;

	assign L1[255:252] = sbox[ in[255:252] ];
	assign L1[251:248] = sbox[ in[251:248] ];
	assign L1[247:244] = sbox[ in[247:244] ];
	assign L1[243:240] = sbox[ in[243:240] ];
	assign L1[239:236] = sbox[ in[239:236] ];
	assign L1[235:232] = sbox[ in[235:232] ];
	assign L1[231:228] = sbox[ in[231:228] ];
	assign L1[227:224] = sbox[ in[227:224] ];
	assign L1[223:220] = sbox[ in[223:220] ];
	assign L1[219:216] = sbox[ in[219:216] ];
	assign L1[215:212] = sbox[ in[215:212] ];
	assign L1[211:208] = sbox[ in[211:208] ];
	assign L1[207:204] = sbox[ in[207:204] ];
	assign L1[203:200] = sbox[ in[203:200] ];
	assign L1[199:196] = sbox[ in[199:196] ];
	assign L1[195:192] = sbox[ in[195:192] ];
	assign L1[191:188] = sbox[ in[191:188] ];
	assign L1[187:184] = sbox[ in[187:184] ];
	assign L1[183:180] = sbox[ in[183:180] ];
	assign L1[179:176] = sbox[ in[179:176] ];
	assign L1[175:172] = sbox[ in[175:172] ];
	assign L1[171:168] = sbox[ in[171:168] ];
	assign L1[167:164] = sbox[ in[167:164] ];
	assign L1[163:160] = sbox[ in[163:160] ];
	assign L1[159:156] = sbox[ in[159:156] ];
	assign L1[155:152] = sbox[ in[155:152] ];
	assign L1[151:148] = sbox[ in[151:148] ];
	assign L1[147:144] = sbox[ in[147:144] ];
	assign L1[143:140] = sbox[ in[143:140] ];
	assign L1[139:136] = sbox[ in[139:136] ];
	assign L1[135:132] = sbox[ in[135:132] ];
	assign L1[131:128] = sbox[ in[131:128] ];
	assign L1[127:124] = sbox[ in[127:124] ];
	assign L1[123:120] = sbox[ in[123:120] ];
	assign L1[119:116] = sbox[ in[119:116] ];
	assign L1[115:112] = sbox[ in[115:112] ];
	assign L1[111:108] = sbox[ in[111:108] ];
	assign L1[107:104] = sbox[ in[107:104] ];
	assign L1[103:100] = sbox[ in[103:100] ];
	assign L1[99:96] = sbox[ in[99:96] ];
	assign L1[95:92] = sbox[ in[95:92] ];
	assign L1[91:88] = sbox[ in[91:88] ];
	assign L1[87:84] = sbox[ in[87:84] ];
	assign L1[83:80] = sbox[ in[83:80] ];
	assign L1[79:76] = sbox[ in[79:76] ];
	assign L1[75:72] = sbox[ in[75:72] ];
	assign L1[71:68] = sbox[ in[71:68] ];
	assign L1[67:64] = sbox[ in[67:64] ];
	assign L1[63:60] = sbox[ in[63:60] ];
	assign L1[59:56] = sbox[ in[59:56] ];
	assign L1[55:52] = sbox[ in[55:52] ];
	assign L1[51:48] = sbox[ in[51:48] ];
	assign L1[47:44] = sbox[ in[47:44] ];
	assign L1[43:40] = sbox[ in[43:40] ];
	assign L1[39:36] = sbox[ in[39:36] ];
	assign L1[35:32] = sbox[ in[35:32] ];
	assign L1[31:28] = sbox[ in[31:28] ];
	assign L1[27:24] = sbox[ in[27:24] ];
	assign L1[23:20] = sbox[ in[23:20] ];
	assign L1[19:16] = sbox[ in[19:16] ];
	assign L1[15:12] = sbox[ in[15:12] ];
	assign L1[11:8] = sbox[ in[11:8] ];
	assign L1[7:4] = sbox[ in[7:4] ];
	assign L1[3:0] = sbox[ in[3:0] ];

	assign out[255:252] = { L1[244]^L1[243], L1[245]^L1[240]^L1[243], L1[246]^L1[241], L1[247]^L1[242] };
	assign out[251:248] = { L1[248]^L1[255]^L1[250], L1[249]^L1[252]^L1[251]^L1[255]^L1[250], L1[250]^L1[253]^L1[248]^L1[251], L1[251]^L1[254]^L1[249] };
	assign out[247:244] = { L1[228]^L1[227], L1[229]^L1[224]^L1[227], L1[230]^L1[225], L1[231]^L1[226] };
	assign out[243:240] = { L1[232]^L1[239]^L1[234], L1[233]^L1[236]^L1[235]^L1[239]^L1[234], L1[234]^L1[237]^L1[232]^L1[235], L1[235]^L1[238]^L1[233] };
	assign out[239:236] = { L1[212]^L1[211], L1[213]^L1[208]^L1[211], L1[214]^L1[209], L1[215]^L1[210] };
	assign out[235:232] = { L1[216]^L1[223]^L1[218], L1[217]^L1[220]^L1[219]^L1[223]^L1[218], L1[218]^L1[221]^L1[216]^L1[219], L1[219]^L1[222]^L1[217] };
	assign out[231:228] = { L1[196]^L1[195], L1[197]^L1[192]^L1[195], L1[198]^L1[193], L1[199]^L1[194] };
	assign out[227:224] = { L1[200]^L1[207]^L1[202], L1[201]^L1[204]^L1[203]^L1[207]^L1[202], L1[202]^L1[205]^L1[200]^L1[203], L1[203]^L1[206]^L1[201] };
	assign out[223:220] = { L1[180]^L1[179], L1[181]^L1[176]^L1[179], L1[182]^L1[177], L1[183]^L1[178] };
	assign out[219:216] = { L1[184]^L1[191]^L1[186], L1[185]^L1[188]^L1[187]^L1[191]^L1[186], L1[186]^L1[189]^L1[184]^L1[187], L1[187]^L1[190]^L1[185] };
	assign out[215:212] = { L1[164]^L1[163], L1[165]^L1[160]^L1[163], L1[166]^L1[161], L1[167]^L1[162] };
	assign out[211:208] = { L1[168]^L1[175]^L1[170], L1[169]^L1[172]^L1[171]^L1[175]^L1[170], L1[170]^L1[173]^L1[168]^L1[171], L1[171]^L1[174]^L1[169] };
	assign out[207:204] = { L1[148]^L1[147], L1[149]^L1[144]^L1[147], L1[150]^L1[145], L1[151]^L1[146] };
	assign out[203:200] = { L1[152]^L1[159]^L1[154], L1[153]^L1[156]^L1[155]^L1[159]^L1[154], L1[154]^L1[157]^L1[152]^L1[155], L1[155]^L1[158]^L1[153] };
	assign out[199:196] = { L1[132]^L1[131], L1[133]^L1[128]^L1[131], L1[134]^L1[129], L1[135]^L1[130] };
	assign out[195:192] = { L1[136]^L1[143]^L1[138], L1[137]^L1[140]^L1[139]^L1[143]^L1[138], L1[138]^L1[141]^L1[136]^L1[139], L1[139]^L1[142]^L1[137] };
	assign out[191:188] = { L1[116]^L1[115], L1[117]^L1[112]^L1[115], L1[118]^L1[113], L1[119]^L1[114] };
	assign out[187:184] = { L1[120]^L1[127]^L1[122], L1[121]^L1[124]^L1[123]^L1[127]^L1[122], L1[122]^L1[125]^L1[120]^L1[123], L1[123]^L1[126]^L1[121] };
	assign out[183:180] = { L1[100]^L1[99], L1[101]^L1[96]^L1[99], L1[102]^L1[97], L1[103]^L1[98] };
	assign out[179:176] = { L1[104]^L1[111]^L1[106], L1[105]^L1[108]^L1[107]^L1[111]^L1[106], L1[106]^L1[109]^L1[104]^L1[107], L1[107]^L1[110]^L1[105] };
	assign out[175:172] = { L1[84]^L1[83], L1[85]^L1[80]^L1[83], L1[86]^L1[81], L1[87]^L1[82] };
	assign out[171:168] = { L1[88]^L1[95]^L1[90], L1[89]^L1[92]^L1[91]^L1[95]^L1[90], L1[90]^L1[93]^L1[88]^L1[91], L1[91]^L1[94]^L1[89] };
	assign out[167:164] = { L1[68]^L1[67], L1[69]^L1[64]^L1[67], L1[70]^L1[65], L1[71]^L1[66] };
	assign out[163:160] = { L1[72]^L1[79]^L1[74], L1[73]^L1[76]^L1[75]^L1[79]^L1[74], L1[74]^L1[77]^L1[72]^L1[75], L1[75]^L1[78]^L1[73] };
	assign out[159:156] = { L1[52]^L1[51], L1[53]^L1[48]^L1[51], L1[54]^L1[49], L1[55]^L1[50] };
	assign out[155:152] = { L1[56]^L1[63]^L1[58], L1[57]^L1[60]^L1[59]^L1[63]^L1[58], L1[58]^L1[61]^L1[56]^L1[59], L1[59]^L1[62]^L1[57] };
	assign out[151:148] = { L1[36]^L1[35], L1[37]^L1[32]^L1[35], L1[38]^L1[33], L1[39]^L1[34] };
	assign out[147:144] = { L1[40]^L1[47]^L1[42], L1[41]^L1[44]^L1[43]^L1[47]^L1[42], L1[42]^L1[45]^L1[40]^L1[43], L1[43]^L1[46]^L1[41] };
	assign out[143:140] = { L1[20]^L1[19], L1[21]^L1[16]^L1[19], L1[22]^L1[17], L1[23]^L1[18] };
	assign out[139:136] = { L1[24]^L1[31]^L1[26], L1[25]^L1[28]^L1[27]^L1[31]^L1[26], L1[26]^L1[29]^L1[24]^L1[27], L1[27]^L1[30]^L1[25] };
	assign out[135:132] = { L1[4]^L1[3], L1[5]^L1[0]^L1[3], L1[6]^L1[1], L1[7]^L1[2] };
	assign out[131:128] = { L1[8]^L1[15]^L1[10], L1[9]^L1[12]^L1[11]^L1[15]^L1[10], L1[10]^L1[13]^L1[8]^L1[11], L1[11]^L1[14]^L1[9] };
	assign out[127:124] = { L1[252]^L1[251], L1[253]^L1[248]^L1[251], L1[254]^L1[249], L1[255]^L1[250] };
	assign out[123:120] = { L1[240]^L1[247]^L1[242], L1[241]^L1[244]^L1[243]^L1[247]^L1[242], L1[242]^L1[245]^L1[240]^L1[243], L1[243]^L1[246]^L1[241] };
	assign out[119:116] = { L1[236]^L1[235], L1[237]^L1[232]^L1[235], L1[238]^L1[233], L1[239]^L1[234] };
	assign out[115:112] = { L1[224]^L1[231]^L1[226], L1[225]^L1[228]^L1[227]^L1[231]^L1[226], L1[226]^L1[229]^L1[224]^L1[227], L1[227]^L1[230]^L1[225] };
	assign out[111:108] = { L1[220]^L1[219], L1[221]^L1[216]^L1[219], L1[222]^L1[217], L1[223]^L1[218] };
	assign out[107:104] = { L1[208]^L1[215]^L1[210], L1[209]^L1[212]^L1[211]^L1[215]^L1[210], L1[210]^L1[213]^L1[208]^L1[211], L1[211]^L1[214]^L1[209] };
	assign out[103:100] = { L1[204]^L1[203], L1[205]^L1[200]^L1[203], L1[206]^L1[201], L1[207]^L1[202] };
	assign out[99:96]   = { L1[192]^L1[199]^L1[194], L1[193]^L1[196]^L1[195]^L1[199]^L1[194], L1[194]^L1[197]^L1[192]^L1[195], L1[195]^L1[198]^L1[193] };
	assign out[95:92]   = { L1[188]^L1[187], L1[189]^L1[184]^L1[187], L1[190]^L1[185], L1[191]^L1[186] };
	assign out[91:88]   = { L1[176]^L1[183]^L1[178], L1[177]^L1[180]^L1[179]^L1[183]^L1[178], L1[178]^L1[181]^L1[176]^L1[179], L1[179]^L1[182]^L1[177] };
	assign out[87:84]   = { L1[172]^L1[171], L1[173]^L1[168]^L1[171], L1[174]^L1[169], L1[175]^L1[170] };
	assign out[83:80]   = { L1[160]^L1[167]^L1[162], L1[161]^L1[164]^L1[163]^L1[167]^L1[162], L1[162]^L1[165]^L1[160]^L1[163], L1[163]^L1[166]^L1[161] };
	assign out[79:76]   = { L1[156]^L1[155], L1[157]^L1[152]^L1[155], L1[158]^L1[153], L1[159]^L1[154] };
	assign out[75:72]   = { L1[144]^L1[151]^L1[146], L1[145]^L1[148]^L1[147]^L1[151]^L1[146], L1[146]^L1[149]^L1[144]^L1[147], L1[147]^L1[150]^L1[145] };
	assign out[71:68]   = { L1[140]^L1[139], L1[141]^L1[136]^L1[139], L1[142]^L1[137], L1[143]^L1[138] };
	assign out[67:64]   = { L1[128]^L1[135]^L1[130], L1[129]^L1[132]^L1[131]^L1[135]^L1[130], L1[130]^L1[133]^L1[128]^L1[131], L1[131]^L1[134]^L1[129] };
	assign out[63:60]   = { L1[124]^L1[123], L1[125]^L1[120]^L1[123], L1[126]^L1[121], L1[127]^L1[122] };
	assign out[59:56]   = { L1[112]^L1[119]^L1[114], L1[113]^L1[116]^L1[115]^L1[119]^L1[114], L1[114]^L1[117]^L1[112]^L1[115], L1[115]^L1[118]^L1[113] };
	assign out[55:52]   = { L1[108]^L1[107], L1[109]^L1[104]^L1[107], L1[110]^L1[105], L1[111]^L1[106] };
	assign out[51:48]   = { L1[96]^L1[103]^L1[98], L1[97]^L1[100]^L1[99]^L1[103]^L1[98], L1[98]^L1[101]^L1[96]^L1[99], L1[99]^L1[102]^L1[97] };
	assign out[47:44]   = { L1[92]^L1[91], L1[93]^L1[88]^L1[91], L1[94]^L1[89], L1[95]^L1[90] };
	assign out[43:40]   = { L1[80]^L1[87]^L1[82], L1[81]^L1[84]^L1[83]^L1[87]^L1[82], L1[82]^L1[85]^L1[80]^L1[83], L1[83]^L1[86]^L1[81] };
	assign out[39:36]   = { L1[76]^L1[75], L1[77]^L1[72]^L1[75], L1[78]^L1[73], L1[79]^L1[74] };
	assign out[35:32]   = { L1[64]^L1[71]^L1[66], L1[65]^L1[68]^L1[67]^L1[71]^L1[66], L1[66]^L1[69]^L1[64]^L1[67], L1[67]^L1[70]^L1[65] };
	assign out[31:28]   = { L1[60]^L1[59], L1[61]^L1[56]^L1[59], L1[62]^L1[57], L1[63]^L1[58] };
	assign out[27:24]   = { L1[48]^L1[55]^L1[50], L1[49]^L1[52]^L1[51]^L1[55]^L1[50], L1[50]^L1[53]^L1[48]^L1[51], L1[51]^L1[54]^L1[49] };
	assign out[23:20]   = { L1[44]^L1[43], L1[45]^L1[40]^L1[43], L1[46]^L1[41], L1[47]^L1[42] };
	assign out[19:16]   = { L1[32]^L1[39]^L1[34], L1[33]^L1[36]^L1[35]^L1[39]^L1[34], L1[34]^L1[37]^L1[32]^L1[35], L1[35]^L1[38]^L1[33] };
	assign out[15:12]   = { L1[28]^L1[27], L1[29]^L1[24]^L1[27], L1[30]^L1[25], L1[31]^L1[26] };
	assign out[11:8]    = { L1[16]^L1[23]^L1[18], L1[17]^L1[20]^L1[19]^L1[23]^L1[18], L1[18]^L1[21]^L1[16]^L1[19], L1[19]^L1[22]^L1[17] };
	assign out[7:4]     = { L1[12]^L1[11], L1[13]^L1[8]^L1[11], L1[14]^L1[9], L1[15]^L1[10] };
	assign out[3:0]     = { L1[0]^L1[7]^L1[2], L1[1]^L1[4]^L1[3]^L1[7]^L1[2], L1[2]^L1[5]^L1[0]^L1[3], L1[3]^L1[6]^L1[1] };

endmodule 

