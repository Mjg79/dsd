module jh_init (
	input [1023:0] in,
	output [1023:0] out
);

	assign out[3:0] = { in[7], in[263], in[519], in[775] };
	assign out[11:8] = { in[6], in[262], in[518], in[774] };
	assign out[19:16] = { in[5], in[261], in[517], in[773] };
	assign out[27:24] = { in[4], in[260], in[516], in[772] };
	assign out[35:32] = { in[3], in[259], in[515], in[771] };
	assign out[43:40] = { in[2], in[258], in[514], in[770] };
	assign out[51:48] = { in[1], in[257], in[513], in[769] };
	assign out[59:56] = { in[0], in[256], in[512], in[768] };
	assign out[67:64] = { in[15], in[271], in[527], in[783] };
	assign out[75:72] = { in[14], in[270], in[526], in[782] };
	assign out[83:80] = { in[13], in[269], in[525], in[781] };
	assign out[91:88] = { in[12], in[268], in[524], in[780] };
	assign out[99:96] = { in[11], in[267], in[523], in[779] };
	assign out[107:104] = { in[10], in[266], in[522], in[778] };
	assign out[115:112] = { in[9], in[265], in[521], in[777] };
	assign out[123:120] = { in[8], in[264], in[520], in[776] };
	assign out[131:128] = { in[23], in[279], in[535], in[791] };
	assign out[139:136] = { in[22], in[278], in[534], in[790] };
	assign out[147:144] = { in[21], in[277], in[533], in[789] };
	assign out[155:152] = { in[20], in[276], in[532], in[788] };
	assign out[163:160] = { in[19], in[275], in[531], in[787] };
	assign out[171:168] = { in[18], in[274], in[530], in[786] };
	assign out[179:176] = { in[17], in[273], in[529], in[785] };
	assign out[187:184] = { in[16], in[272], in[528], in[784] };
	assign out[195:192] = { in[31], in[287], in[543], in[799] };
	assign out[203:200] = { in[30], in[286], in[542], in[798] };
	assign out[211:208] = { in[29], in[285], in[541], in[797] };
	assign out[219:216] = { in[28], in[284], in[540], in[796] };
	assign out[227:224] = { in[27], in[283], in[539], in[795] };
	assign out[235:232] = { in[26], in[282], in[538], in[794] };
	assign out[243:240] = { in[25], in[281], in[537], in[793] };
	assign out[251:248] = { in[24], in[280], in[536], in[792] };
	assign out[259:256] = { in[39], in[295], in[551], in[807] };
	assign out[267:264] = { in[38], in[294], in[550], in[806] };
	assign out[275:272] = { in[37], in[293], in[549], in[805] };
	assign out[283:280] = { in[36], in[292], in[548], in[804] };
	assign out[291:288] = { in[35], in[291], in[547], in[803] };
	assign out[299:296] = { in[34], in[290], in[546], in[802] };
	assign out[307:304] = { in[33], in[289], in[545], in[801] };
	assign out[315:312] = { in[32], in[288], in[544], in[800] };
	assign out[323:320] = { in[47], in[303], in[559], in[815] };
	assign out[331:328] = { in[46], in[302], in[558], in[814] };
	assign out[339:336] = { in[45], in[301], in[557], in[813] };
	assign out[347:344] = { in[44], in[300], in[556], in[812] };
	assign out[355:352] = { in[43], in[299], in[555], in[811] };
	assign out[363:360] = { in[42], in[298], in[554], in[810] };
	assign out[371:368] = { in[41], in[297], in[553], in[809] };
	assign out[379:376] = { in[40], in[296], in[552], in[808] };
	assign out[387:384] = { in[55], in[311], in[567], in[823] };
	assign out[395:392] = { in[54], in[310], in[566], in[822] };
	assign out[403:400] = { in[53], in[309], in[565], in[821] };
	assign out[411:408] = { in[52], in[308], in[564], in[820] };
	assign out[419:416] = { in[51], in[307], in[563], in[819] };
	assign out[427:424] = { in[50], in[306], in[562], in[818] };
	assign out[435:432] = { in[49], in[305], in[561], in[817] };
	assign out[443:440] = { in[48], in[304], in[560], in[816] };
	assign out[451:448] = { in[63], in[319], in[575], in[831] };
	assign out[459:456] = { in[62], in[318], in[574], in[830] };
	assign out[467:464] = { in[61], in[317], in[573], in[829] };
	assign out[475:472] = { in[60], in[316], in[572], in[828] };
	assign out[483:480] = { in[59], in[315], in[571], in[827] };
	assign out[491:488] = { in[58], in[314], in[570], in[826] };
	assign out[499:496] = { in[57], in[313], in[569], in[825] };
	assign out[507:504] = { in[56], in[312], in[568], in[824] };
	assign out[515:512] = { in[71], in[327], in[583], in[839] };
	assign out[523:520] = { in[70], in[326], in[582], in[838] };
	assign out[531:528] = { in[69], in[325], in[581], in[837] };
	assign out[539:536] = { in[68], in[324], in[580], in[836] };
	assign out[547:544] = { in[67], in[323], in[579], in[835] };
	assign out[555:552] = { in[66], in[322], in[578], in[834] };
	assign out[563:560] = { in[65], in[321], in[577], in[833] };
	assign out[571:568] = { in[64], in[320], in[576], in[832] };
	assign out[579:576] = { in[79], in[335], in[591], in[847] };
	assign out[587:584] = { in[78], in[334], in[590], in[846] };
	assign out[595:592] = { in[77], in[333], in[589], in[845] };
	assign out[603:600] = { in[76], in[332], in[588], in[844] };
	assign out[611:608] = { in[75], in[331], in[587], in[843] };
	assign out[619:616] = { in[74], in[330], in[586], in[842] };
	assign out[627:624] = { in[73], in[329], in[585], in[841] };
	assign out[635:632] = { in[72], in[328], in[584], in[840] };
	assign out[643:640] = { in[87], in[343], in[599], in[855] };
	assign out[651:648] = { in[86], in[342], in[598], in[854] };
	assign out[659:656] = { in[85], in[341], in[597], in[853] };
	assign out[667:664] = { in[84], in[340], in[596], in[852] };
	assign out[675:672] = { in[83], in[339], in[595], in[851] };
	assign out[683:680] = { in[82], in[338], in[594], in[850] };
	assign out[691:688] = { in[81], in[337], in[593], in[849] };
	assign out[699:696] = { in[80], in[336], in[592], in[848] };
	assign out[707:704] = { in[95], in[351], in[607], in[863] };
	assign out[715:712] = { in[94], in[350], in[606], in[862] };
	assign out[723:720] = { in[93], in[349], in[605], in[861] };
	assign out[731:728] = { in[92], in[348], in[604], in[860] };
	assign out[739:736] = { in[91], in[347], in[603], in[859] };
	assign out[747:744] = { in[90], in[346], in[602], in[858] };
	assign out[755:752] = { in[89], in[345], in[601], in[857] };
	assign out[763:760] = { in[88], in[344], in[600], in[856] };
	assign out[771:768] = { in[103], in[359], in[615], in[871] };
	assign out[779:776] = { in[102], in[358], in[614], in[870] };
	assign out[787:784] = { in[101], in[357], in[613], in[869] };
	assign out[795:792] = { in[100], in[356], in[612], in[868] };
	assign out[803:800] = { in[99], in[355], in[611], in[867] };
	assign out[811:808] = { in[98], in[354], in[610], in[866] };
	assign out[819:816] = { in[97], in[353], in[609], in[865] };
	assign out[827:824] = { in[96], in[352], in[608], in[864] };
	assign out[835:832] = { in[111], in[367], in[623], in[879] };
	assign out[843:840] = { in[110], in[366], in[622], in[878] };
	assign out[851:848] = { in[109], in[365], in[621], in[877] };
	assign out[859:856] = { in[108], in[364], in[620], in[876] };
	assign out[867:864] = { in[107], in[363], in[619], in[875] };
	assign out[875:872] = { in[106], in[362], in[618], in[874] };
	assign out[883:880] = { in[105], in[361], in[617], in[873] };
	assign out[891:888] = { in[104], in[360], in[616], in[872] };
	assign out[899:896] = { in[119], in[375], in[631], in[887] };
	assign out[907:904] = { in[118], in[374], in[630], in[886] };
	assign out[915:912] = { in[117], in[373], in[629], in[885] };
	assign out[923:920] = { in[116], in[372], in[628], in[884] };
	assign out[931:928] = { in[115], in[371], in[627], in[883] };
	assign out[939:936] = { in[114], in[370], in[626], in[882] };
	assign out[947:944] = { in[113], in[369], in[625], in[881] };
	assign out[955:952] = { in[112], in[368], in[624], in[880] };
	assign out[963:960] = { in[127], in[383], in[639], in[895] };
	assign out[971:968] = { in[126], in[382], in[638], in[894] };
	assign out[979:976] = { in[125], in[381], in[637], in[893] };
	assign out[987:984] = { in[124], in[380], in[636], in[892] };
	assign out[995:992] = { in[123], in[379], in[635], in[891] };
	assign out[1003:1000] = { in[122], in[378], in[634], in[890] };
	assign out[1011:1008] = { in[121], in[377], in[633], in[889] };
	assign out[1019:1016] = { in[120], in[376], in[632], in[888] };
	assign out[7:4] = { in[135], in[391], in[647], in[903] };
	assign out[15:12] = { in[134], in[390], in[646], in[902] };
	assign out[23:20] = { in[133], in[389], in[645], in[901] };
	assign out[31:28] = { in[132], in[388], in[644], in[900] };
	assign out[39:36] = { in[131], in[387], in[643], in[899] };
	assign out[47:44] = { in[130], in[386], in[642], in[898] };
	assign out[55:52] = { in[129], in[385], in[641], in[897] };
	assign out[63:60] = { in[128], in[384], in[640], in[896] };
	assign out[71:68] = { in[143], in[399], in[655], in[911] };
	assign out[79:76] = { in[142], in[398], in[654], in[910] };
	assign out[87:84] = { in[141], in[397], in[653], in[909] };
	assign out[95:92] = { in[140], in[396], in[652], in[908] };
	assign out[103:100] = { in[139], in[395], in[651], in[907] };
	assign out[111:108] = { in[138], in[394], in[650], in[906] };
	assign out[119:116] = { in[137], in[393], in[649], in[905] };
	assign out[127:124] = { in[136], in[392], in[648], in[904] };
	assign out[135:132] = { in[151], in[407], in[663], in[919] };
	assign out[143:140] = { in[150], in[406], in[662], in[918] };
	assign out[151:148] = { in[149], in[405], in[661], in[917] };
	assign out[159:156] = { in[148], in[404], in[660], in[916] };
	assign out[167:164] = { in[147], in[403], in[659], in[915] };
	assign out[175:172] = { in[146], in[402], in[658], in[914] };
	assign out[183:180] = { in[145], in[401], in[657], in[913] };
	assign out[191:188] = { in[144], in[400], in[656], in[912] };
	assign out[199:196] = { in[159], in[415], in[671], in[927] };
	assign out[207:204] = { in[158], in[414], in[670], in[926] };
	assign out[215:212] = { in[157], in[413], in[669], in[925] };
	assign out[223:220] = { in[156], in[412], in[668], in[924] };
	assign out[231:228] = { in[155], in[411], in[667], in[923] };
	assign out[239:236] = { in[154], in[410], in[666], in[922] };
	assign out[247:244] = { in[153], in[409], in[665], in[921] };
	assign out[255:252] = { in[152], in[408], in[664], in[920] };
	assign out[263:260] = { in[167], in[423], in[679], in[935] };
	assign out[271:268] = { in[166], in[422], in[678], in[934] };
	assign out[279:276] = { in[165], in[421], in[677], in[933] };
	assign out[287:284] = { in[164], in[420], in[676], in[932] };
	assign out[295:292] = { in[163], in[419], in[675], in[931] };
	assign out[303:300] = { in[162], in[418], in[674], in[930] };
	assign out[311:308] = { in[161], in[417], in[673], in[929] };
	assign out[319:316] = { in[160], in[416], in[672], in[928] };
	assign out[327:324] = { in[175], in[431], in[687], in[943] };
	assign out[335:332] = { in[174], in[430], in[686], in[942] };
	assign out[343:340] = { in[173], in[429], in[685], in[941] };
	assign out[351:348] = { in[172], in[428], in[684], in[940] };
	assign out[359:356] = { in[171], in[427], in[683], in[939] };
	assign out[367:364] = { in[170], in[426], in[682], in[938] };
	assign out[375:372] = { in[169], in[425], in[681], in[937] };
	assign out[383:380] = { in[168], in[424], in[680], in[936] };
	assign out[391:388] = { in[183], in[439], in[695], in[951] };
	assign out[399:396] = { in[182], in[438], in[694], in[950] };
	assign out[407:404] = { in[181], in[437], in[693], in[949] };
	assign out[415:412] = { in[180], in[436], in[692], in[948] };
	assign out[423:420] = { in[179], in[435], in[691], in[947] };
	assign out[431:428] = { in[178], in[434], in[690], in[946] };
	assign out[439:436] = { in[177], in[433], in[689], in[945] };
	assign out[447:444] = { in[176], in[432], in[688], in[944] };
	assign out[455:452] = { in[191], in[447], in[703], in[959] };
	assign out[463:460] = { in[190], in[446], in[702], in[958] };
	assign out[471:468] = { in[189], in[445], in[701], in[957] };
	assign out[479:476] = { in[188], in[444], in[700], in[956] };
	assign out[487:484] = { in[187], in[443], in[699], in[955] };
	assign out[495:492] = { in[186], in[442], in[698], in[954] };
	assign out[503:500] = { in[185], in[441], in[697], in[953] };
	assign out[511:508] = { in[184], in[440], in[696], in[952] };
	assign out[519:516] = { in[199], in[455], in[711], in[967] };
	assign out[527:524] = { in[198], in[454], in[710], in[966] };
	assign out[535:532] = { in[197], in[453], in[709], in[965] };
	assign out[543:540] = { in[196], in[452], in[708], in[964] };
	assign out[551:548] = { in[195], in[451], in[707], in[963] };
	assign out[559:556] = { in[194], in[450], in[706], in[962] };
	assign out[567:564] = { in[193], in[449], in[705], in[961] };
	assign out[575:572] = { in[192], in[448], in[704], in[960] };
	assign out[583:580] = { in[207], in[463], in[719], in[975] };
	assign out[591:588] = { in[206], in[462], in[718], in[974] };
	assign out[599:596] = { in[205], in[461], in[717], in[973] };
	assign out[607:604] = { in[204], in[460], in[716], in[972] };
	assign out[615:612] = { in[203], in[459], in[715], in[971] };
	assign out[623:620] = { in[202], in[458], in[714], in[970] };
	assign out[631:628] = { in[201], in[457], in[713], in[969] };
	assign out[639:636] = { in[200], in[456], in[712], in[968] };
	assign out[647:644] = { in[215], in[471], in[727], in[983] };
	assign out[655:652] = { in[214], in[470], in[726], in[982] };
	assign out[663:660] = { in[213], in[469], in[725], in[981] };
	assign out[671:668] = { in[212], in[468], in[724], in[980] };
	assign out[679:676] = { in[211], in[467], in[723], in[979] };
	assign out[687:684] = { in[210], in[466], in[722], in[978] };
	assign out[695:692] = { in[209], in[465], in[721], in[977] };
	assign out[703:700] = { in[208], in[464], in[720], in[976] };
	assign out[711:708] = { in[223], in[479], in[735], in[991] };
	assign out[719:716] = { in[222], in[478], in[734], in[990] };
	assign out[727:724] = { in[221], in[477], in[733], in[989] };
	assign out[735:732] = { in[220], in[476], in[732], in[988] };
	assign out[743:740] = { in[219], in[475], in[731], in[987] };
	assign out[751:748] = { in[218], in[474], in[730], in[986] };
	assign out[759:756] = { in[217], in[473], in[729], in[985] };
	assign out[767:764] = { in[216], in[472], in[728], in[984] };
	assign out[775:772] = { in[231], in[487], in[743], in[999] };
	assign out[783:780] = { in[230], in[486], in[742], in[998] };
	assign out[791:788] = { in[229], in[485], in[741], in[997] };
	assign out[799:796] = { in[228], in[484], in[740], in[996] };
	assign out[807:804] = { in[227], in[483], in[739], in[995] };
	assign out[815:812] = { in[226], in[482], in[738], in[994] };
	assign out[823:820] = { in[225], in[481], in[737], in[993] };
	assign out[831:828] = { in[224], in[480], in[736], in[992] };
	assign out[839:836] = { in[239], in[495], in[751], in[1007] };
	assign out[847:844] = { in[238], in[494], in[750], in[1006] };
	assign out[855:852] = { in[237], in[493], in[749], in[1005] };
	assign out[863:860] = { in[236], in[492], in[748], in[1004] };
	assign out[871:868] = { in[235], in[491], in[747], in[1003] };
	assign out[879:876] = { in[234], in[490], in[746], in[1002] };
	assign out[887:884] = { in[233], in[489], in[745], in[1001] };
	assign out[895:892] = { in[232], in[488], in[744], in[1000] };
	assign out[903:900] = { in[247], in[503], in[759], in[1015] };
	assign out[911:908] = { in[246], in[502], in[758], in[1014] };
	assign out[919:916] = { in[245], in[501], in[757], in[1013] };
	assign out[927:924] = { in[244], in[500], in[756], in[1012] };
	assign out[935:932] = { in[243], in[499], in[755], in[1011] };
	assign out[943:940] = { in[242], in[498], in[754], in[1010] };
	assign out[951:948] = { in[241], in[497], in[753], in[1009] };
	assign out[959:956] = { in[240], in[496], in[752], in[1008] };
	assign out[967:964] = { in[255], in[511], in[767], in[1023] };
	assign out[975:972] = { in[254], in[510], in[766], in[1022] };
	assign out[983:980] = { in[253], in[509], in[765], in[1021] };
	assign out[991:988] = { in[252], in[508], in[764], in[1020] };
	assign out[999:996] = { in[251], in[507], in[763], in[1019] };
	assign out[1007:1004] = { in[250], in[506], in[762], in[1018] };
	assign out[1015:1012] = { in[249], in[505], in[761], in[1017] };
	assign out[1023:1020] = { in[248], in[504], in[760], in[1016] };
	
endmodule

