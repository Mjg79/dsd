module jh_round_a (
	input [1023:0] state_in,
	input [255:0] round_in,
	output [1023:0] out
);         

	wire [3:0] sbox [0:31] = { 4'h9,4'h0,4'h4,4'hb,4'hd,4'hc,4'h3,4'hf,4'h1,4'ha,4'h2,4'h6,4'h7,4'h5,4'h8,4'he,4'h3,4'hc,4'h6,4'hd,4'h5,4'h7,4'h1,4'h9,4'hf,4'h2,4'h0,4'h4,4'hb,4'ha,4'he,4'h8 };
	
	wire [1023:0] L1;

	assign L1[1023:1020] = sbox[ { round_in[255], state_in[1023:1020] } ];
	assign L1[1019:1016] = sbox[ { round_in[254], state_in[1019:1016] } ];
	assign L1[1015:1012] = sbox[ { round_in[253], state_in[1015:1012] } ];
	assign L1[1011:1008] = sbox[ { round_in[252], state_in[1011:1008] } ];
	assign L1[1007:1004] = sbox[ { round_in[251], state_in[1007:1004] } ];
	assign L1[1003:1000] = sbox[ { round_in[250], state_in[1003:1000] } ];
	assign L1[999:996] = sbox[ { round_in[249], state_in[999:996] } ];
	assign L1[995:992] = sbox[ { round_in[248], state_in[995:992] } ];
	assign L1[991:988] = sbox[ { round_in[247], state_in[991:988] } ];
	assign L1[987:984] = sbox[ { round_in[246], state_in[987:984] } ];
	assign L1[983:980] = sbox[ { round_in[245], state_in[983:980] } ];
	assign L1[979:976] = sbox[ { round_in[244], state_in[979:976] } ];
	assign L1[975:972] = sbox[ { round_in[243], state_in[975:972] } ];
	assign L1[971:968] = sbox[ { round_in[242], state_in[971:968] } ];
	assign L1[967:964] = sbox[ { round_in[241], state_in[967:964] } ];
	assign L1[963:960] = sbox[ { round_in[240], state_in[963:960] } ];
	assign L1[959:956] = sbox[ { round_in[239], state_in[959:956] } ];
	assign L1[955:952] = sbox[ { round_in[238], state_in[955:952] } ];
	assign L1[951:948] = sbox[ { round_in[237], state_in[951:948] } ];
	assign L1[947:944] = sbox[ { round_in[236], state_in[947:944] } ];
	assign L1[943:940] = sbox[ { round_in[235], state_in[943:940] } ];
	assign L1[939:936] = sbox[ { round_in[234], state_in[939:936] } ];
	assign L1[935:932] = sbox[ { round_in[233], state_in[935:932] } ];
	assign L1[931:928] = sbox[ { round_in[232], state_in[931:928] } ];
	assign L1[927:924] = sbox[ { round_in[231], state_in[927:924] } ];
	assign L1[923:920] = sbox[ { round_in[230], state_in[923:920] } ];
	assign L1[919:916] = sbox[ { round_in[229], state_in[919:916] } ];
	assign L1[915:912] = sbox[ { round_in[228], state_in[915:912] } ];
	assign L1[911:908] = sbox[ { round_in[227], state_in[911:908] } ];
	assign L1[907:904] = sbox[ { round_in[226], state_in[907:904] } ];
	assign L1[903:900] = sbox[ { round_in[225], state_in[903:900] } ];
	assign L1[899:896] = sbox[ { round_in[224], state_in[899:896] } ];
	assign L1[895:892] = sbox[ { round_in[223], state_in[895:892] } ];
	assign L1[891:888] = sbox[ { round_in[222], state_in[891:888] } ];
	assign L1[887:884] = sbox[ { round_in[221], state_in[887:884] } ];
	assign L1[883:880] = sbox[ { round_in[220], state_in[883:880] } ];
	assign L1[879:876] = sbox[ { round_in[219], state_in[879:876] } ];
	assign L1[875:872] = sbox[ { round_in[218], state_in[875:872] } ];
	assign L1[871:868] = sbox[ { round_in[217], state_in[871:868] } ];
	assign L1[867:864] = sbox[ { round_in[216], state_in[867:864] } ];
	assign L1[863:860] = sbox[ { round_in[215], state_in[863:860] } ];
	assign L1[859:856] = sbox[ { round_in[214], state_in[859:856] } ];
	assign L1[855:852] = sbox[ { round_in[213], state_in[855:852] } ];
	assign L1[851:848] = sbox[ { round_in[212], state_in[851:848] } ];
	assign L1[847:844] = sbox[ { round_in[211], state_in[847:844] } ];
	assign L1[843:840] = sbox[ { round_in[210], state_in[843:840] } ];
	assign L1[839:836] = sbox[ { round_in[209], state_in[839:836] } ];
	assign L1[835:832] = sbox[ { round_in[208], state_in[835:832] } ];
	assign L1[831:828] = sbox[ { round_in[207], state_in[831:828] } ];
	assign L1[827:824] = sbox[ { round_in[206], state_in[827:824] } ];
	assign L1[823:820] = sbox[ { round_in[205], state_in[823:820] } ];
	assign L1[819:816] = sbox[ { round_in[204], state_in[819:816] } ];
	assign L1[815:812] = sbox[ { round_in[203], state_in[815:812] } ];
	assign L1[811:808] = sbox[ { round_in[202], state_in[811:808] } ];
	assign L1[807:804] = sbox[ { round_in[201], state_in[807:804] } ];
	assign L1[803:800] = sbox[ { round_in[200], state_in[803:800] } ];
	assign L1[799:796] = sbox[ { round_in[199], state_in[799:796] } ];
	assign L1[795:792] = sbox[ { round_in[198], state_in[795:792] } ];
	assign L1[791:788] = sbox[ { round_in[197], state_in[791:788] } ];
	assign L1[787:784] = sbox[ { round_in[196], state_in[787:784] } ];
	assign L1[783:780] = sbox[ { round_in[195], state_in[783:780] } ];
	assign L1[779:776] = sbox[ { round_in[194], state_in[779:776] } ];
	assign L1[775:772] = sbox[ { round_in[193], state_in[775:772] } ];
	assign L1[771:768] = sbox[ { round_in[192], state_in[771:768] } ];
	assign L1[767:764] = sbox[ { round_in[191], state_in[767:764] } ];
	assign L1[763:760] = sbox[ { round_in[190], state_in[763:760] } ];
	assign L1[759:756] = sbox[ { round_in[189], state_in[759:756] } ];
	assign L1[755:752] = sbox[ { round_in[188], state_in[755:752] } ];
	assign L1[751:748] = sbox[ { round_in[187], state_in[751:748] } ];
	assign L1[747:744] = sbox[ { round_in[186], state_in[747:744] } ];
	assign L1[743:740] = sbox[ { round_in[185], state_in[743:740] } ];
	assign L1[739:736] = sbox[ { round_in[184], state_in[739:736] } ];
	assign L1[735:732] = sbox[ { round_in[183], state_in[735:732] } ];
	assign L1[731:728] = sbox[ { round_in[182], state_in[731:728] } ];
	assign L1[727:724] = sbox[ { round_in[181], state_in[727:724] } ];
	assign L1[723:720] = sbox[ { round_in[180], state_in[723:720] } ];
	assign L1[719:716] = sbox[ { round_in[179], state_in[719:716] } ];
	assign L1[715:712] = sbox[ { round_in[178], state_in[715:712] } ];
	assign L1[711:708] = sbox[ { round_in[177], state_in[711:708] } ];
	assign L1[707:704] = sbox[ { round_in[176], state_in[707:704] } ];
	assign L1[703:700] = sbox[ { round_in[175], state_in[703:700] } ];
	assign L1[699:696] = sbox[ { round_in[174], state_in[699:696] } ];
	assign L1[695:692] = sbox[ { round_in[173], state_in[695:692] } ];
	assign L1[691:688] = sbox[ { round_in[172], state_in[691:688] } ];
	assign L1[687:684] = sbox[ { round_in[171], state_in[687:684] } ];
	assign L1[683:680] = sbox[ { round_in[170], state_in[683:680] } ];
	assign L1[679:676] = sbox[ { round_in[169], state_in[679:676] } ];
	assign L1[675:672] = sbox[ { round_in[168], state_in[675:672] } ];
	assign L1[671:668] = sbox[ { round_in[167], state_in[671:668] } ];
	assign L1[667:664] = sbox[ { round_in[166], state_in[667:664] } ];
	assign L1[663:660] = sbox[ { round_in[165], state_in[663:660] } ];
	assign L1[659:656] = sbox[ { round_in[164], state_in[659:656] } ];
	assign L1[655:652] = sbox[ { round_in[163], state_in[655:652] } ];
	assign L1[651:648] = sbox[ { round_in[162], state_in[651:648] } ];
	assign L1[647:644] = sbox[ { round_in[161], state_in[647:644] } ];
	assign L1[643:640] = sbox[ { round_in[160], state_in[643:640] } ];
	assign L1[639:636] = sbox[ { round_in[159], state_in[639:636] } ];
	assign L1[635:632] = sbox[ { round_in[158], state_in[635:632] } ];
	assign L1[631:628] = sbox[ { round_in[157], state_in[631:628] } ];
	assign L1[627:624] = sbox[ { round_in[156], state_in[627:624] } ];
	assign L1[623:620] = sbox[ { round_in[155], state_in[623:620] } ];
	assign L1[619:616] = sbox[ { round_in[154], state_in[619:616] } ];
	assign L1[615:612] = sbox[ { round_in[153], state_in[615:612] } ];
	assign L1[611:608] = sbox[ { round_in[152], state_in[611:608] } ];
	assign L1[607:604] = sbox[ { round_in[151], state_in[607:604] } ];
	assign L1[603:600] = sbox[ { round_in[150], state_in[603:600] } ];
	assign L1[599:596] = sbox[ { round_in[149], state_in[599:596] } ];
	assign L1[595:592] = sbox[ { round_in[148], state_in[595:592] } ];
	assign L1[591:588] = sbox[ { round_in[147], state_in[591:588] } ];
	assign L1[587:584] = sbox[ { round_in[146], state_in[587:584] } ];
	assign L1[583:580] = sbox[ { round_in[145], state_in[583:580] } ];
	assign L1[579:576] = sbox[ { round_in[144], state_in[579:576] } ];
	assign L1[575:572] = sbox[ { round_in[143], state_in[575:572] } ];
	assign L1[571:568] = sbox[ { round_in[142], state_in[571:568] } ];
	assign L1[567:564] = sbox[ { round_in[141], state_in[567:564] } ];
	assign L1[563:560] = sbox[ { round_in[140], state_in[563:560] } ];
	assign L1[559:556] = sbox[ { round_in[139], state_in[559:556] } ];
	assign L1[555:552] = sbox[ { round_in[138], state_in[555:552] } ];
	assign L1[551:548] = sbox[ { round_in[137], state_in[551:548] } ];
	assign L1[547:544] = sbox[ { round_in[136], state_in[547:544] } ];
	assign L1[543:540] = sbox[ { round_in[135], state_in[543:540] } ];
	assign L1[539:536] = sbox[ { round_in[134], state_in[539:536] } ];
	assign L1[535:532] = sbox[ { round_in[133], state_in[535:532] } ];
	assign L1[531:528] = sbox[ { round_in[132], state_in[531:528] } ];
	assign L1[527:524] = sbox[ { round_in[131], state_in[527:524] } ];
	assign L1[523:520] = sbox[ { round_in[130], state_in[523:520] } ];
	assign L1[519:516] = sbox[ { round_in[129], state_in[519:516] } ];
	assign L1[515:512] = sbox[ { round_in[128], state_in[515:512] } ];
	assign L1[511:508] = sbox[ { round_in[127], state_in[511:508] } ];
	assign L1[507:504] = sbox[ { round_in[126], state_in[507:504] } ];
	assign L1[503:500] = sbox[ { round_in[125], state_in[503:500] } ];
	assign L1[499:496] = sbox[ { round_in[124], state_in[499:496] } ];
	assign L1[495:492] = sbox[ { round_in[123], state_in[495:492] } ];
	assign L1[491:488] = sbox[ { round_in[122], state_in[491:488] } ];
	assign L1[487:484] = sbox[ { round_in[121], state_in[487:484] } ];
	assign L1[483:480] = sbox[ { round_in[120], state_in[483:480] } ];
	assign L1[479:476] = sbox[ { round_in[119], state_in[479:476] } ];
	assign L1[475:472] = sbox[ { round_in[118], state_in[475:472] } ];
	assign L1[471:468] = sbox[ { round_in[117], state_in[471:468] } ];
	assign L1[467:464] = sbox[ { round_in[116], state_in[467:464] } ];
	assign L1[463:460] = sbox[ { round_in[115], state_in[463:460] } ];
	assign L1[459:456] = sbox[ { round_in[114], state_in[459:456] } ];
	assign L1[455:452] = sbox[ { round_in[113], state_in[455:452] } ];
	assign L1[451:448] = sbox[ { round_in[112], state_in[451:448] } ];
	assign L1[447:444] = sbox[ { round_in[111], state_in[447:444] } ];
	assign L1[443:440] = sbox[ { round_in[110], state_in[443:440] } ];
	assign L1[439:436] = sbox[ { round_in[109], state_in[439:436] } ];
	assign L1[435:432] = sbox[ { round_in[108], state_in[435:432] } ];
	assign L1[431:428] = sbox[ { round_in[107], state_in[431:428] } ];
	assign L1[427:424] = sbox[ { round_in[106], state_in[427:424] } ];
	assign L1[423:420] = sbox[ { round_in[105], state_in[423:420] } ];
	assign L1[419:416] = sbox[ { round_in[104], state_in[419:416] } ];
	assign L1[415:412] = sbox[ { round_in[103], state_in[415:412] } ];
	assign L1[411:408] = sbox[ { round_in[102], state_in[411:408] } ];
	assign L1[407:404] = sbox[ { round_in[101], state_in[407:404] } ];
	assign L1[403:400] = sbox[ { round_in[100], state_in[403:400] } ];
	assign L1[399:396] = sbox[ { round_in[99], state_in[399:396] } ];
	assign L1[395:392] = sbox[ { round_in[98], state_in[395:392] } ];
	assign L1[391:388] = sbox[ { round_in[97], state_in[391:388] } ];
	assign L1[387:384] = sbox[ { round_in[96], state_in[387:384] } ];
	assign L1[383:380] = sbox[ { round_in[95], state_in[383:380] } ];
	assign L1[379:376] = sbox[ { round_in[94], state_in[379:376] } ];
	assign L1[375:372] = sbox[ { round_in[93], state_in[375:372] } ];
	assign L1[371:368] = sbox[ { round_in[92], state_in[371:368] } ];
	assign L1[367:364] = sbox[ { round_in[91], state_in[367:364] } ];
	assign L1[363:360] = sbox[ { round_in[90], state_in[363:360] } ];
	assign L1[359:356] = sbox[ { round_in[89], state_in[359:356] } ];
	assign L1[355:352] = sbox[ { round_in[88], state_in[355:352] } ];
	assign L1[351:348] = sbox[ { round_in[87], state_in[351:348] } ];
	assign L1[347:344] = sbox[ { round_in[86], state_in[347:344] } ];
	assign L1[343:340] = sbox[ { round_in[85], state_in[343:340] } ];
	assign L1[339:336] = sbox[ { round_in[84], state_in[339:336] } ];
	assign L1[335:332] = sbox[ { round_in[83], state_in[335:332] } ];
	assign L1[331:328] = sbox[ { round_in[82], state_in[331:328] } ];
	assign L1[327:324] = sbox[ { round_in[81], state_in[327:324] } ];
	assign L1[323:320] = sbox[ { round_in[80], state_in[323:320] } ];
	assign L1[319:316] = sbox[ { round_in[79], state_in[319:316] } ];
	assign L1[315:312] = sbox[ { round_in[78], state_in[315:312] } ];
	assign L1[311:308] = sbox[ { round_in[77], state_in[311:308] } ];
	assign L1[307:304] = sbox[ { round_in[76], state_in[307:304] } ];
	assign L1[303:300] = sbox[ { round_in[75], state_in[303:300] } ];
	assign L1[299:296] = sbox[ { round_in[74], state_in[299:296] } ];
	assign L1[295:292] = sbox[ { round_in[73], state_in[295:292] } ];
	assign L1[291:288] = sbox[ { round_in[72], state_in[291:288] } ];
	assign L1[287:284] = sbox[ { round_in[71], state_in[287:284] } ];
	assign L1[283:280] = sbox[ { round_in[70], state_in[283:280] } ];
	assign L1[279:276] = sbox[ { round_in[69], state_in[279:276] } ];
	assign L1[275:272] = sbox[ { round_in[68], state_in[275:272] } ];
	assign L1[271:268] = sbox[ { round_in[67], state_in[271:268] } ];
	assign L1[267:264] = sbox[ { round_in[66], state_in[267:264] } ];
	assign L1[263:260] = sbox[ { round_in[65], state_in[263:260] } ];
	assign L1[259:256] = sbox[ { round_in[64], state_in[259:256] } ];
	assign L1[255:252] = sbox[ { round_in[63], state_in[255:252] } ];
	assign L1[251:248] = sbox[ { round_in[62], state_in[251:248] } ];
	assign L1[247:244] = sbox[ { round_in[61], state_in[247:244] } ];
	assign L1[243:240] = sbox[ { round_in[60], state_in[243:240] } ];
	assign L1[239:236] = sbox[ { round_in[59], state_in[239:236] } ];
	assign L1[235:232] = sbox[ { round_in[58], state_in[235:232] } ];
	assign L1[231:228] = sbox[ { round_in[57], state_in[231:228] } ];
	assign L1[227:224] = sbox[ { round_in[56], state_in[227:224] } ];
	assign L1[223:220] = sbox[ { round_in[55], state_in[223:220] } ];
	assign L1[219:216] = sbox[ { round_in[54], state_in[219:216] } ];
	assign L1[215:212] = sbox[ { round_in[53], state_in[215:212] } ];
	assign L1[211:208] = sbox[ { round_in[52], state_in[211:208] } ];
	assign L1[207:204] = sbox[ { round_in[51], state_in[207:204] } ];
	assign L1[203:200] = sbox[ { round_in[50], state_in[203:200] } ];
	assign L1[199:196] = sbox[ { round_in[49], state_in[199:196] } ];
	assign L1[195:192] = sbox[ { round_in[48], state_in[195:192] } ];
	assign L1[191:188] = sbox[ { round_in[47], state_in[191:188] } ];
	assign L1[187:184] = sbox[ { round_in[46], state_in[187:184] } ];
	assign L1[183:180] = sbox[ { round_in[45], state_in[183:180] } ];
	assign L1[179:176] = sbox[ { round_in[44], state_in[179:176] } ];
	assign L1[175:172] = sbox[ { round_in[43], state_in[175:172] } ];
	assign L1[171:168] = sbox[ { round_in[42], state_in[171:168] } ];
	assign L1[167:164] = sbox[ { round_in[41], state_in[167:164] } ];
	assign L1[163:160] = sbox[ { round_in[40], state_in[163:160] } ];
	assign L1[159:156] = sbox[ { round_in[39], state_in[159:156] } ];
	assign L1[155:152] = sbox[ { round_in[38], state_in[155:152] } ];
	assign L1[151:148] = sbox[ { round_in[37], state_in[151:148] } ];
	assign L1[147:144] = sbox[ { round_in[36], state_in[147:144] } ];
	assign L1[143:140] = sbox[ { round_in[35], state_in[143:140] } ];
	assign L1[139:136] = sbox[ { round_in[34], state_in[139:136] } ];
	assign L1[135:132] = sbox[ { round_in[33], state_in[135:132] } ];
	assign L1[131:128] = sbox[ { round_in[32], state_in[131:128] } ];
	assign L1[127:124] = sbox[ { round_in[31], state_in[127:124] } ];
	assign L1[123:120] = sbox[ { round_in[30], state_in[123:120] } ];
	assign L1[119:116] = sbox[ { round_in[29], state_in[119:116] } ];
	assign L1[115:112] = sbox[ { round_in[28], state_in[115:112] } ];
	assign L1[111:108] = sbox[ { round_in[27], state_in[111:108] } ];
	assign L1[107:104] = sbox[ { round_in[26], state_in[107:104] } ];
	assign L1[103:100] = sbox[ { round_in[25], state_in[103:100] } ];
	assign L1[99:96] = sbox[ { round_in[24], state_in[99:96] } ];
	assign L1[95:92] = sbox[ { round_in[23], state_in[95:92] } ];
	assign L1[91:88] = sbox[ { round_in[22], state_in[91:88] } ];
	assign L1[87:84] = sbox[ { round_in[21], state_in[87:84] } ];
	assign L1[83:80] = sbox[ { round_in[20], state_in[83:80] } ];
	assign L1[79:76] = sbox[ { round_in[19], state_in[79:76] } ];
	assign L1[75:72] = sbox[ { round_in[18], state_in[75:72] } ];
	assign L1[71:68] = sbox[ { round_in[17], state_in[71:68] } ];
	assign L1[67:64] = sbox[ { round_in[16], state_in[67:64] } ];
	assign L1[63:60] = sbox[ { round_in[15], state_in[63:60] } ];
	assign L1[59:56] = sbox[ { round_in[14], state_in[59:56] } ];
	assign L1[55:52] = sbox[ { round_in[13], state_in[55:52] } ];
	assign L1[51:48] = sbox[ { round_in[12], state_in[51:48] } ];
	assign L1[47:44] = sbox[ { round_in[11], state_in[47:44] } ];
	assign L1[43:40] = sbox[ { round_in[10], state_in[43:40] } ];
	assign L1[39:36] = sbox[ { round_in[9], state_in[39:36] } ];
	assign L1[35:32] = sbox[ { round_in[8], state_in[35:32] } ];
	assign L1[31:28] = sbox[ { round_in[7], state_in[31:28] } ];
	assign L1[27:24] = sbox[ { round_in[6], state_in[27:24] } ];
	assign L1[23:20] = sbox[ { round_in[5], state_in[23:20] } ];
	assign L1[19:16] = sbox[ { round_in[4], state_in[19:16] } ];
	assign L1[15:12] = sbox[ { round_in[3], state_in[15:12] } ];
	assign L1[11:8] = sbox[ { round_in[2], state_in[11:8] } ];
	assign L1[7:4] = sbox[ { round_in[1], state_in[7:4] } ];
	assign L1[3:0] = sbox[ { round_in[0], state_in[3:0] } ];

	assign out[1023:1020] = { L1[1015]^L1[1010], L1[1014]^L1[1009], L1[1013]^L1[1008]^L1[1011], L1[1012]^L1[1011] };
	assign out[1019:1016] = { L1[1019]^L1[1022]^L1[1017], L1[1018]^L1[1021]^L1[1016]^L1[1019], L1[1017]^L1[1020]^L1[1019]^L1[1023]^L1[1018], L1[1016]^L1[1023]^L1[1018] };
	assign out[1015:1012] = { L1[999]^L1[994], L1[998]^L1[993], L1[997]^L1[992]^L1[995], L1[996]^L1[995] };
	assign out[1011:1008] = { L1[1003]^L1[1006]^L1[1001], L1[1002]^L1[1005]^L1[1000]^L1[1003], L1[1001]^L1[1004]^L1[1003]^L1[1007]^L1[1002], L1[1000]^L1[1007]^L1[1002] };
	assign out[1007:1004] = { L1[983]^L1[978], L1[982]^L1[977], L1[981]^L1[976]^L1[979], L1[980]^L1[979] };
	assign out[1003:1000] = { L1[987]^L1[990]^L1[985], L1[986]^L1[989]^L1[984]^L1[987], L1[985]^L1[988]^L1[987]^L1[991]^L1[986], L1[984]^L1[991]^L1[986] };
	assign out[999:996]   = { L1[967]^L1[962], L1[966]^L1[961], L1[965]^L1[960]^L1[963], L1[964]^L1[963] };
	assign out[995:992]   = { L1[971]^L1[974]^L1[969], L1[970]^L1[973]^L1[968]^L1[971], L1[969]^L1[972]^L1[971]^L1[975]^L1[970], L1[968]^L1[975]^L1[970] };
	assign out[991:988]   = { L1[951]^L1[946], L1[950]^L1[945], L1[949]^L1[944]^L1[947], L1[948]^L1[947] };
	assign out[987:984]   = { L1[955]^L1[958]^L1[953], L1[954]^L1[957]^L1[952]^L1[955], L1[953]^L1[956]^L1[955]^L1[959]^L1[954], L1[952]^L1[959]^L1[954] };
	assign out[983:980]   = { L1[935]^L1[930], L1[934]^L1[929], L1[933]^L1[928]^L1[931], L1[932]^L1[931] };
	assign out[979:976]   = { L1[939]^L1[942]^L1[937], L1[938]^L1[941]^L1[936]^L1[939], L1[937]^L1[940]^L1[939]^L1[943]^L1[938], L1[936]^L1[943]^L1[938] };
	assign out[975:972]   = { L1[919]^L1[914], L1[918]^L1[913], L1[917]^L1[912]^L1[915], L1[916]^L1[915] };
	assign out[971:968]   = { L1[923]^L1[926]^L1[921], L1[922]^L1[925]^L1[920]^L1[923], L1[921]^L1[924]^L1[923]^L1[927]^L1[922], L1[920]^L1[927]^L1[922] };
	assign out[967:964]   = { L1[903]^L1[898], L1[902]^L1[897], L1[901]^L1[896]^L1[899], L1[900]^L1[899] };
	assign out[963:960]   = { L1[907]^L1[910]^L1[905], L1[906]^L1[909]^L1[904]^L1[907], L1[905]^L1[908]^L1[907]^L1[911]^L1[906], L1[904]^L1[911]^L1[906] };
	assign out[959:956]   = { L1[887]^L1[882], L1[886]^L1[881], L1[885]^L1[880]^L1[883], L1[884]^L1[883] };
	assign out[955:952]   = { L1[891]^L1[894]^L1[889], L1[890]^L1[893]^L1[888]^L1[891], L1[889]^L1[892]^L1[891]^L1[895]^L1[890], L1[888]^L1[895]^L1[890] };
	assign out[951:948]   = { L1[871]^L1[866], L1[870]^L1[865], L1[869]^L1[864]^L1[867], L1[868]^L1[867] };
	assign out[947:944]   = { L1[875]^L1[878]^L1[873], L1[874]^L1[877]^L1[872]^L1[875], L1[873]^L1[876]^L1[875]^L1[879]^L1[874], L1[872]^L1[879]^L1[874] };
	assign out[943:940]   = { L1[855]^L1[850], L1[854]^L1[849], L1[853]^L1[848]^L1[851], L1[852]^L1[851] };
	assign out[939:936]   = { L1[859]^L1[862]^L1[857], L1[858]^L1[861]^L1[856]^L1[859], L1[857]^L1[860]^L1[859]^L1[863]^L1[858], L1[856]^L1[863]^L1[858] };
	assign out[935:932]   = { L1[839]^L1[834], L1[838]^L1[833], L1[837]^L1[832]^L1[835], L1[836]^L1[835] };
	assign out[931:928]   = { L1[843]^L1[846]^L1[841], L1[842]^L1[845]^L1[840]^L1[843], L1[841]^L1[844]^L1[843]^L1[847]^L1[842], L1[840]^L1[847]^L1[842] };
	assign out[927:924]   = { L1[823]^L1[818], L1[822]^L1[817], L1[821]^L1[816]^L1[819], L1[820]^L1[819] };
	assign out[923:920]   = { L1[827]^L1[830]^L1[825], L1[826]^L1[829]^L1[824]^L1[827], L1[825]^L1[828]^L1[827]^L1[831]^L1[826], L1[824]^L1[831]^L1[826] };
	assign out[919:916]   = { L1[807]^L1[802], L1[806]^L1[801], L1[805]^L1[800]^L1[803], L1[804]^L1[803] };
	assign out[915:912]   = { L1[811]^L1[814]^L1[809], L1[810]^L1[813]^L1[808]^L1[811], L1[809]^L1[812]^L1[811]^L1[815]^L1[810], L1[808]^L1[815]^L1[810] };
	assign out[911:908]   = { L1[791]^L1[786], L1[790]^L1[785], L1[789]^L1[784]^L1[787], L1[788]^L1[787] };
	assign out[907:904]   = { L1[795]^L1[798]^L1[793], L1[794]^L1[797]^L1[792]^L1[795], L1[793]^L1[796]^L1[795]^L1[799]^L1[794], L1[792]^L1[799]^L1[794] };
	assign out[903:900]   = { L1[775]^L1[770], L1[774]^L1[769], L1[773]^L1[768]^L1[771], L1[772]^L1[771] };
	assign out[899:896]   = { L1[779]^L1[782]^L1[777], L1[778]^L1[781]^L1[776]^L1[779], L1[777]^L1[780]^L1[779]^L1[783]^L1[778], L1[776]^L1[783]^L1[778] };
	assign out[895:892]   = { L1[759]^L1[754], L1[758]^L1[753], L1[757]^L1[752]^L1[755], L1[756]^L1[755] };
	assign out[891:888]   = { L1[763]^L1[766]^L1[761], L1[762]^L1[765]^L1[760]^L1[763], L1[761]^L1[764]^L1[763]^L1[767]^L1[762], L1[760]^L1[767]^L1[762] };
	assign out[887:884]   = { L1[743]^L1[738], L1[742]^L1[737], L1[741]^L1[736]^L1[739], L1[740]^L1[739] };
	assign out[883:880]   = { L1[747]^L1[750]^L1[745], L1[746]^L1[749]^L1[744]^L1[747], L1[745]^L1[748]^L1[747]^L1[751]^L1[746], L1[744]^L1[751]^L1[746] };
	assign out[879:876]   = { L1[727]^L1[722], L1[726]^L1[721], L1[725]^L1[720]^L1[723], L1[724]^L1[723] };
	assign out[875:872]   = { L1[731]^L1[734]^L1[729], L1[730]^L1[733]^L1[728]^L1[731], L1[729]^L1[732]^L1[731]^L1[735]^L1[730], L1[728]^L1[735]^L1[730] };
	assign out[871:868]   = { L1[711]^L1[706], L1[710]^L1[705], L1[709]^L1[704]^L1[707], L1[708]^L1[707] };
	assign out[867:864]   = { L1[715]^L1[718]^L1[713], L1[714]^L1[717]^L1[712]^L1[715], L1[713]^L1[716]^L1[715]^L1[719]^L1[714], L1[712]^L1[719]^L1[714] };
	assign out[863:860]   = { L1[695]^L1[690], L1[694]^L1[689], L1[693]^L1[688]^L1[691], L1[692]^L1[691] };
	assign out[859:856]   = { L1[699]^L1[702]^L1[697], L1[698]^L1[701]^L1[696]^L1[699], L1[697]^L1[700]^L1[699]^L1[703]^L1[698], L1[696]^L1[703]^L1[698] };
	assign out[855:852]   = { L1[679]^L1[674], L1[678]^L1[673], L1[677]^L1[672]^L1[675], L1[676]^L1[675] };
	assign out[851:848]   = { L1[683]^L1[686]^L1[681], L1[682]^L1[685]^L1[680]^L1[683], L1[681]^L1[684]^L1[683]^L1[687]^L1[682], L1[680]^L1[687]^L1[682] };
	assign out[847:844]   = { L1[663]^L1[658], L1[662]^L1[657], L1[661]^L1[656]^L1[659], L1[660]^L1[659] };
	assign out[843:840]   = { L1[667]^L1[670]^L1[665], L1[666]^L1[669]^L1[664]^L1[667], L1[665]^L1[668]^L1[667]^L1[671]^L1[666], L1[664]^L1[671]^L1[666] };
	assign out[839:836]   = { L1[647]^L1[642], L1[646]^L1[641], L1[645]^L1[640]^L1[643], L1[644]^L1[643] };
	assign out[835:832]   = { L1[651]^L1[654]^L1[649], L1[650]^L1[653]^L1[648]^L1[651], L1[649]^L1[652]^L1[651]^L1[655]^L1[650], L1[648]^L1[655]^L1[650] };
	assign out[831:828]   = { L1[631]^L1[626], L1[630]^L1[625], L1[629]^L1[624]^L1[627], L1[628]^L1[627] };
	assign out[827:824]   = { L1[635]^L1[638]^L1[633], L1[634]^L1[637]^L1[632]^L1[635], L1[633]^L1[636]^L1[635]^L1[639]^L1[634], L1[632]^L1[639]^L1[634] };
	assign out[823:820]   = { L1[615]^L1[610], L1[614]^L1[609], L1[613]^L1[608]^L1[611], L1[612]^L1[611] };
	assign out[819:816]   = { L1[619]^L1[622]^L1[617], L1[618]^L1[621]^L1[616]^L1[619], L1[617]^L1[620]^L1[619]^L1[623]^L1[618], L1[616]^L1[623]^L1[618] };
	assign out[815:812]   = { L1[599]^L1[594], L1[598]^L1[593], L1[597]^L1[592]^L1[595], L1[596]^L1[595] };
	assign out[811:808]   = { L1[603]^L1[606]^L1[601], L1[602]^L1[605]^L1[600]^L1[603], L1[601]^L1[604]^L1[603]^L1[607]^L1[602], L1[600]^L1[607]^L1[602] };
	assign out[807:804]   = { L1[583]^L1[578], L1[582]^L1[577], L1[581]^L1[576]^L1[579], L1[580]^L1[579] };
	assign out[803:800]   = { L1[587]^L1[590]^L1[585], L1[586]^L1[589]^L1[584]^L1[587], L1[585]^L1[588]^L1[587]^L1[591]^L1[586], L1[584]^L1[591]^L1[586] };
	assign out[799:796]   = { L1[567]^L1[562], L1[566]^L1[561], L1[565]^L1[560]^L1[563], L1[564]^L1[563] };
	assign out[795:792]   = { L1[571]^L1[574]^L1[569], L1[570]^L1[573]^L1[568]^L1[571], L1[569]^L1[572]^L1[571]^L1[575]^L1[570], L1[568]^L1[575]^L1[570] };
	assign out[791:788]   = { L1[551]^L1[546], L1[550]^L1[545], L1[549]^L1[544]^L1[547], L1[548]^L1[547] };
	assign out[787:784]   = { L1[555]^L1[558]^L1[553], L1[554]^L1[557]^L1[552]^L1[555], L1[553]^L1[556]^L1[555]^L1[559]^L1[554], L1[552]^L1[559]^L1[554] };
	assign out[783:780]   = { L1[535]^L1[530], L1[534]^L1[529], L1[533]^L1[528]^L1[531], L1[532]^L1[531] };
	assign out[779:776]   = { L1[539]^L1[542]^L1[537], L1[538]^L1[541]^L1[536]^L1[539], L1[537]^L1[540]^L1[539]^L1[543]^L1[538], L1[536]^L1[543]^L1[538] };
	assign out[775:772]   = { L1[519]^L1[514], L1[518]^L1[513], L1[517]^L1[512]^L1[515], L1[516]^L1[515] };
	assign out[771:768]   = { L1[523]^L1[526]^L1[521], L1[522]^L1[525]^L1[520]^L1[523], L1[521]^L1[524]^L1[523]^L1[527]^L1[522], L1[520]^L1[527]^L1[522] };
	assign out[767:764]   = { L1[503]^L1[498], L1[502]^L1[497], L1[501]^L1[496]^L1[499], L1[500]^L1[499] };
	assign out[763:760]   = { L1[507]^L1[510]^L1[505], L1[506]^L1[509]^L1[504]^L1[507], L1[505]^L1[508]^L1[507]^L1[511]^L1[506], L1[504]^L1[511]^L1[506] };
	assign out[759:756]   = { L1[487]^L1[482], L1[486]^L1[481], L1[485]^L1[480]^L1[483], L1[484]^L1[483] };
	assign out[755:752]   = { L1[491]^L1[494]^L1[489], L1[490]^L1[493]^L1[488]^L1[491], L1[489]^L1[492]^L1[491]^L1[495]^L1[490], L1[488]^L1[495]^L1[490] };
	assign out[751:748]   = { L1[471]^L1[466], L1[470]^L1[465], L1[469]^L1[464]^L1[467], L1[468]^L1[467] };
	assign out[747:744]   = { L1[475]^L1[478]^L1[473], L1[474]^L1[477]^L1[472]^L1[475], L1[473]^L1[476]^L1[475]^L1[479]^L1[474], L1[472]^L1[479]^L1[474] };
	assign out[743:740]   = { L1[455]^L1[450], L1[454]^L1[449], L1[453]^L1[448]^L1[451], L1[452]^L1[451] };
	assign out[739:736]   = { L1[459]^L1[462]^L1[457], L1[458]^L1[461]^L1[456]^L1[459], L1[457]^L1[460]^L1[459]^L1[463]^L1[458], L1[456]^L1[463]^L1[458] };
	assign out[735:732]   = { L1[439]^L1[434], L1[438]^L1[433], L1[437]^L1[432]^L1[435], L1[436]^L1[435] };
	assign out[731:728]   = { L1[443]^L1[446]^L1[441], L1[442]^L1[445]^L1[440]^L1[443], L1[441]^L1[444]^L1[443]^L1[447]^L1[442], L1[440]^L1[447]^L1[442] };
	assign out[727:724]   = { L1[423]^L1[418], L1[422]^L1[417], L1[421]^L1[416]^L1[419], L1[420]^L1[419] };
	assign out[723:720]   = { L1[427]^L1[430]^L1[425], L1[426]^L1[429]^L1[424]^L1[427], L1[425]^L1[428]^L1[427]^L1[431]^L1[426], L1[424]^L1[431]^L1[426] };
	assign out[719:716]   = { L1[407]^L1[402], L1[406]^L1[401], L1[405]^L1[400]^L1[403], L1[404]^L1[403] };
	assign out[715:712]   = { L1[411]^L1[414]^L1[409], L1[410]^L1[413]^L1[408]^L1[411], L1[409]^L1[412]^L1[411]^L1[415]^L1[410], L1[408]^L1[415]^L1[410] };
	assign out[711:708]   = { L1[391]^L1[386], L1[390]^L1[385], L1[389]^L1[384]^L1[387], L1[388]^L1[387] };
	assign out[707:704]   = { L1[395]^L1[398]^L1[393], L1[394]^L1[397]^L1[392]^L1[395], L1[393]^L1[396]^L1[395]^L1[399]^L1[394], L1[392]^L1[399]^L1[394] };
	assign out[703:700]   = { L1[375]^L1[370], L1[374]^L1[369], L1[373]^L1[368]^L1[371], L1[372]^L1[371] };
	assign out[699:696]   = { L1[379]^L1[382]^L1[377], L1[378]^L1[381]^L1[376]^L1[379], L1[377]^L1[380]^L1[379]^L1[383]^L1[378], L1[376]^L1[383]^L1[378] };
	assign out[695:692]   = { L1[359]^L1[354], L1[358]^L1[353], L1[357]^L1[352]^L1[355], L1[356]^L1[355] };
	assign out[691:688]   = { L1[363]^L1[366]^L1[361], L1[362]^L1[365]^L1[360]^L1[363], L1[361]^L1[364]^L1[363]^L1[367]^L1[362], L1[360]^L1[367]^L1[362] };
	assign out[687:684]   = { L1[343]^L1[338], L1[342]^L1[337], L1[341]^L1[336]^L1[339], L1[340]^L1[339] };
	assign out[683:680]   = { L1[347]^L1[350]^L1[345], L1[346]^L1[349]^L1[344]^L1[347], L1[345]^L1[348]^L1[347]^L1[351]^L1[346], L1[344]^L1[351]^L1[346] };
	assign out[679:676]   = { L1[327]^L1[322], L1[326]^L1[321], L1[325]^L1[320]^L1[323], L1[324]^L1[323] };
	assign out[675:672]   = { L1[331]^L1[334]^L1[329], L1[330]^L1[333]^L1[328]^L1[331], L1[329]^L1[332]^L1[331]^L1[335]^L1[330], L1[328]^L1[335]^L1[330] };
	assign out[671:668]   = { L1[311]^L1[306], L1[310]^L1[305], L1[309]^L1[304]^L1[307], L1[308]^L1[307] };
	assign out[667:664]   = { L1[315]^L1[318]^L1[313], L1[314]^L1[317]^L1[312]^L1[315], L1[313]^L1[316]^L1[315]^L1[319]^L1[314], L1[312]^L1[319]^L1[314] };
	assign out[663:660]   = { L1[295]^L1[290], L1[294]^L1[289], L1[293]^L1[288]^L1[291], L1[292]^L1[291] };
	assign out[659:656]   = { L1[299]^L1[302]^L1[297], L1[298]^L1[301]^L1[296]^L1[299], L1[297]^L1[300]^L1[299]^L1[303]^L1[298], L1[296]^L1[303]^L1[298] };
	assign out[655:652]   = { L1[279]^L1[274], L1[278]^L1[273], L1[277]^L1[272]^L1[275], L1[276]^L1[275] };
	assign out[651:648]   = { L1[283]^L1[286]^L1[281], L1[282]^L1[285]^L1[280]^L1[283], L1[281]^L1[284]^L1[283]^L1[287]^L1[282], L1[280]^L1[287]^L1[282] };
	assign out[647:644]   = { L1[263]^L1[258], L1[262]^L1[257], L1[261]^L1[256]^L1[259], L1[260]^L1[259] };
	assign out[643:640]   = { L1[267]^L1[270]^L1[265], L1[266]^L1[269]^L1[264]^L1[267], L1[265]^L1[268]^L1[267]^L1[271]^L1[266], L1[264]^L1[271]^L1[266] };
	assign out[639:636]   = { L1[247]^L1[242], L1[246]^L1[241], L1[245]^L1[240]^L1[243], L1[244]^L1[243] };
	assign out[635:632]   = { L1[251]^L1[254]^L1[249], L1[250]^L1[253]^L1[248]^L1[251], L1[249]^L1[252]^L1[251]^L1[255]^L1[250], L1[248]^L1[255]^L1[250] };
	assign out[631:628]   = { L1[231]^L1[226], L1[230]^L1[225], L1[229]^L1[224]^L1[227], L1[228]^L1[227] };
	assign out[627:624]   = { L1[235]^L1[238]^L1[233], L1[234]^L1[237]^L1[232]^L1[235], L1[233]^L1[236]^L1[235]^L1[239]^L1[234], L1[232]^L1[239]^L1[234] };
	assign out[623:620]   = { L1[215]^L1[210], L1[214]^L1[209], L1[213]^L1[208]^L1[211], L1[212]^L1[211] };
	assign out[619:616]   = { L1[219]^L1[222]^L1[217], L1[218]^L1[221]^L1[216]^L1[219], L1[217]^L1[220]^L1[219]^L1[223]^L1[218], L1[216]^L1[223]^L1[218] };
	assign out[615:612]   = { L1[199]^L1[194], L1[198]^L1[193], L1[197]^L1[192]^L1[195], L1[196]^L1[195] };
	assign out[611:608]   = { L1[203]^L1[206]^L1[201], L1[202]^L1[205]^L1[200]^L1[203], L1[201]^L1[204]^L1[203]^L1[207]^L1[202], L1[200]^L1[207]^L1[202] };
	assign out[607:604]   = { L1[183]^L1[178], L1[182]^L1[177], L1[181]^L1[176]^L1[179], L1[180]^L1[179] };
	assign out[603:600]   = { L1[187]^L1[190]^L1[185], L1[186]^L1[189]^L1[184]^L1[187], L1[185]^L1[188]^L1[187]^L1[191]^L1[186], L1[184]^L1[191]^L1[186] };
	assign out[599:596]   = { L1[167]^L1[162], L1[166]^L1[161], L1[165]^L1[160]^L1[163], L1[164]^L1[163] };
	assign out[595:592]   = { L1[171]^L1[174]^L1[169], L1[170]^L1[173]^L1[168]^L1[171], L1[169]^L1[172]^L1[171]^L1[175]^L1[170], L1[168]^L1[175]^L1[170] };
	assign out[591:588]   = { L1[151]^L1[146], L1[150]^L1[145], L1[149]^L1[144]^L1[147], L1[148]^L1[147] };
	assign out[587:584]   = { L1[155]^L1[158]^L1[153], L1[154]^L1[157]^L1[152]^L1[155], L1[153]^L1[156]^L1[155]^L1[159]^L1[154], L1[152]^L1[159]^L1[154] };
	assign out[583:580]   = { L1[135]^L1[130], L1[134]^L1[129], L1[133]^L1[128]^L1[131], L1[132]^L1[131] };
	assign out[579:576]   = { L1[139]^L1[142]^L1[137], L1[138]^L1[141]^L1[136]^L1[139], L1[137]^L1[140]^L1[139]^L1[143]^L1[138], L1[136]^L1[143]^L1[138] };
	assign out[575:572]   = { L1[119]^L1[114], L1[118]^L1[113], L1[117]^L1[112]^L1[115], L1[116]^L1[115] };
	assign out[571:568]   = { L1[123]^L1[126]^L1[121], L1[122]^L1[125]^L1[120]^L1[123], L1[121]^L1[124]^L1[123]^L1[127]^L1[122], L1[120]^L1[127]^L1[122] };
	assign out[567:564]   = { L1[103]^L1[98], L1[102]^L1[97], L1[101]^L1[96]^L1[99], L1[100]^L1[99] };
	assign out[563:560]   = { L1[107]^L1[110]^L1[105], L1[106]^L1[109]^L1[104]^L1[107], L1[105]^L1[108]^L1[107]^L1[111]^L1[106], L1[104]^L1[111]^L1[106] };
	assign out[559:556]   = { L1[87]^L1[82], L1[86]^L1[81], L1[85]^L1[80]^L1[83], L1[84]^L1[83] };
	assign out[555:552]   = { L1[91]^L1[94]^L1[89], L1[90]^L1[93]^L1[88]^L1[91], L1[89]^L1[92]^L1[91]^L1[95]^L1[90], L1[88]^L1[95]^L1[90] };
	assign out[551:548]   = { L1[71]^L1[66], L1[70]^L1[65], L1[69]^L1[64]^L1[67], L1[68]^L1[67] };
	assign out[547:544]   = { L1[75]^L1[78]^L1[73], L1[74]^L1[77]^L1[72]^L1[75], L1[73]^L1[76]^L1[75]^L1[79]^L1[74], L1[72]^L1[79]^L1[74] };
	assign out[543:540]   = { L1[55]^L1[50], L1[54]^L1[49], L1[53]^L1[48]^L1[51], L1[52]^L1[51] };
	assign out[539:536]   = { L1[59]^L1[62]^L1[57], L1[58]^L1[61]^L1[56]^L1[59], L1[57]^L1[60]^L1[59]^L1[63]^L1[58], L1[56]^L1[63]^L1[58] };
	assign out[535:532]   = { L1[39]^L1[34], L1[38]^L1[33], L1[37]^L1[32]^L1[35], L1[36]^L1[35] };
	assign out[531:528]   = { L1[43]^L1[46]^L1[41], L1[42]^L1[45]^L1[40]^L1[43], L1[41]^L1[44]^L1[43]^L1[47]^L1[42], L1[40]^L1[47]^L1[42] };
	assign out[527:524]   = { L1[23]^L1[18], L1[22]^L1[17], L1[21]^L1[16]^L1[19], L1[20]^L1[19] };
	assign out[523:520]   = { L1[27]^L1[30]^L1[25], L1[26]^L1[29]^L1[24]^L1[27], L1[25]^L1[28]^L1[27]^L1[31]^L1[26], L1[24]^L1[31]^L1[26] };
	assign out[519:516]   = { L1[7]^L1[2], L1[6]^L1[1], L1[5]^L1[0]^L1[3], L1[4]^L1[3] };
	assign out[515:512]   = { L1[11]^L1[14]^L1[9], L1[10]^L1[13]^L1[8]^L1[11], L1[9]^L1[12]^L1[11]^L1[15]^L1[10], L1[8]^L1[15]^L1[10] };
	assign out[511:508]   = { L1[1023]^L1[1018], L1[1022]^L1[1017], L1[1021]^L1[1016]^L1[1019], L1[1020]^L1[1019] };
	assign out[507:504]   = { L1[1011]^L1[1014]^L1[1009], L1[1010]^L1[1013]^L1[1008]^L1[1011], L1[1009]^L1[1012]^L1[1011]^L1[1015]^L1[1010], L1[1008]^L1[1015]^L1[1010] };
	assign out[503:500]   = { L1[1007]^L1[1002], L1[1006]^L1[1001], L1[1005]^L1[1000]^L1[1003], L1[1004]^L1[1003] };
	assign out[499:496]   = { L1[995]^L1[998]^L1[993], L1[994]^L1[997]^L1[992]^L1[995], L1[993]^L1[996]^L1[995]^L1[999]^L1[994], L1[992]^L1[999]^L1[994] };
	assign out[495:492]   = { L1[991]^L1[986], L1[990]^L1[985], L1[989]^L1[984]^L1[987], L1[988]^L1[987] };
	assign out[491:488]   = { L1[979]^L1[982]^L1[977], L1[978]^L1[981]^L1[976]^L1[979], L1[977]^L1[980]^L1[979]^L1[983]^L1[978], L1[976]^L1[983]^L1[978] };
	assign out[487:484]   = { L1[975]^L1[970], L1[974]^L1[969], L1[973]^L1[968]^L1[971], L1[972]^L1[971] };
	assign out[483:480]   = { L1[963]^L1[966]^L1[961], L1[962]^L1[965]^L1[960]^L1[963], L1[961]^L1[964]^L1[963]^L1[967]^L1[962], L1[960]^L1[967]^L1[962] };
	assign out[479:476]   = { L1[959]^L1[954], L1[958]^L1[953], L1[957]^L1[952]^L1[955], L1[956]^L1[955] };
	assign out[475:472]   = { L1[947]^L1[950]^L1[945], L1[946]^L1[949]^L1[944]^L1[947], L1[945]^L1[948]^L1[947]^L1[951]^L1[946], L1[944]^L1[951]^L1[946] };
	assign out[471:468]   = { L1[943]^L1[938], L1[942]^L1[937], L1[941]^L1[936]^L1[939], L1[940]^L1[939] };
	assign out[467:464]   = { L1[931]^L1[934]^L1[929], L1[930]^L1[933]^L1[928]^L1[931], L1[929]^L1[932]^L1[931]^L1[935]^L1[930], L1[928]^L1[935]^L1[930] };
	assign out[463:460]   = { L1[927]^L1[922], L1[926]^L1[921], L1[925]^L1[920]^L1[923], L1[924]^L1[923] };
	assign out[459:456]   = { L1[915]^L1[918]^L1[913], L1[914]^L1[917]^L1[912]^L1[915], L1[913]^L1[916]^L1[915]^L1[919]^L1[914], L1[912]^L1[919]^L1[914] };
	assign out[455:452]   = { L1[911]^L1[906], L1[910]^L1[905], L1[909]^L1[904]^L1[907], L1[908]^L1[907] };
	assign out[451:448]   = { L1[899]^L1[902]^L1[897], L1[898]^L1[901]^L1[896]^L1[899], L1[897]^L1[900]^L1[899]^L1[903]^L1[898], L1[896]^L1[903]^L1[898] };
	assign out[447:444]   = { L1[895]^L1[890], L1[894]^L1[889], L1[893]^L1[888]^L1[891], L1[892]^L1[891] };
	assign out[443:440]   = { L1[883]^L1[886]^L1[881], L1[882]^L1[885]^L1[880]^L1[883], L1[881]^L1[884]^L1[883]^L1[887]^L1[882], L1[880]^L1[887]^L1[882] };
	assign out[439:436]   = { L1[879]^L1[874], L1[878]^L1[873], L1[877]^L1[872]^L1[875], L1[876]^L1[875] };
	assign out[435:432]   = { L1[867]^L1[870]^L1[865], L1[866]^L1[869]^L1[864]^L1[867], L1[865]^L1[868]^L1[867]^L1[871]^L1[866], L1[864]^L1[871]^L1[866] };
	assign out[431:428]   = { L1[863]^L1[858], L1[862]^L1[857], L1[861]^L1[856]^L1[859], L1[860]^L1[859] };
	assign out[427:424]   = { L1[851]^L1[854]^L1[849], L1[850]^L1[853]^L1[848]^L1[851], L1[849]^L1[852]^L1[851]^L1[855]^L1[850], L1[848]^L1[855]^L1[850] };
	assign out[423:420]   = { L1[847]^L1[842], L1[846]^L1[841], L1[845]^L1[840]^L1[843], L1[844]^L1[843] };
	assign out[419:416]   = { L1[835]^L1[838]^L1[833], L1[834]^L1[837]^L1[832]^L1[835], L1[833]^L1[836]^L1[835]^L1[839]^L1[834], L1[832]^L1[839]^L1[834] };
	assign out[415:412]   = { L1[831]^L1[826], L1[830]^L1[825], L1[829]^L1[824]^L1[827], L1[828]^L1[827] };
	assign out[411:408]   = { L1[819]^L1[822]^L1[817], L1[818]^L1[821]^L1[816]^L1[819], L1[817]^L1[820]^L1[819]^L1[823]^L1[818], L1[816]^L1[823]^L1[818] };
	assign out[407:404]   = { L1[815]^L1[810], L1[814]^L1[809], L1[813]^L1[808]^L1[811], L1[812]^L1[811] };
	assign out[403:400]   = { L1[803]^L1[806]^L1[801], L1[802]^L1[805]^L1[800]^L1[803], L1[801]^L1[804]^L1[803]^L1[807]^L1[802], L1[800]^L1[807]^L1[802] };
	assign out[399:396]   = { L1[799]^L1[794], L1[798]^L1[793], L1[797]^L1[792]^L1[795], L1[796]^L1[795] };
	assign out[395:392]   = { L1[787]^L1[790]^L1[785], L1[786]^L1[789]^L1[784]^L1[787], L1[785]^L1[788]^L1[787]^L1[791]^L1[786], L1[784]^L1[791]^L1[786] };
	assign out[391:388]   = { L1[783]^L1[778], L1[782]^L1[777], L1[781]^L1[776]^L1[779], L1[780]^L1[779] };
	assign out[387:384]   = { L1[771]^L1[774]^L1[769], L1[770]^L1[773]^L1[768]^L1[771], L1[769]^L1[772]^L1[771]^L1[775]^L1[770], L1[768]^L1[775]^L1[770] };
	assign out[383:380]   = { L1[767]^L1[762], L1[766]^L1[761], L1[765]^L1[760]^L1[763], L1[764]^L1[763] };
	assign out[379:376]   = { L1[755]^L1[758]^L1[753], L1[754]^L1[757]^L1[752]^L1[755], L1[753]^L1[756]^L1[755]^L1[759]^L1[754], L1[752]^L1[759]^L1[754] };
	assign out[375:372]   = { L1[751]^L1[746], L1[750]^L1[745], L1[749]^L1[744]^L1[747], L1[748]^L1[747] };
	assign out[371:368]   = { L1[739]^L1[742]^L1[737], L1[738]^L1[741]^L1[736]^L1[739], L1[737]^L1[740]^L1[739]^L1[743]^L1[738], L1[736]^L1[743]^L1[738] };
	assign out[367:364]   = { L1[735]^L1[730], L1[734]^L1[729], L1[733]^L1[728]^L1[731], L1[732]^L1[731] };
	assign out[363:360]   = { L1[723]^L1[726]^L1[721], L1[722]^L1[725]^L1[720]^L1[723], L1[721]^L1[724]^L1[723]^L1[727]^L1[722], L1[720]^L1[727]^L1[722] };
	assign out[359:356]   = { L1[719]^L1[714], L1[718]^L1[713], L1[717]^L1[712]^L1[715], L1[716]^L1[715] };
	assign out[355:352]   = { L1[707]^L1[710]^L1[705], L1[706]^L1[709]^L1[704]^L1[707], L1[705]^L1[708]^L1[707]^L1[711]^L1[706], L1[704]^L1[711]^L1[706] };
	assign out[351:348]   = { L1[703]^L1[698], L1[702]^L1[697], L1[701]^L1[696]^L1[699], L1[700]^L1[699] };
	assign out[347:344]   = { L1[691]^L1[694]^L1[689], L1[690]^L1[693]^L1[688]^L1[691], L1[689]^L1[692]^L1[691]^L1[695]^L1[690], L1[688]^L1[695]^L1[690] };
	assign out[343:340]   = { L1[687]^L1[682], L1[686]^L1[681], L1[685]^L1[680]^L1[683], L1[684]^L1[683] };
	assign out[339:336]   = { L1[675]^L1[678]^L1[673], L1[674]^L1[677]^L1[672]^L1[675], L1[673]^L1[676]^L1[675]^L1[679]^L1[674], L1[672]^L1[679]^L1[674] };
	assign out[335:332]   = { L1[671]^L1[666], L1[670]^L1[665], L1[669]^L1[664]^L1[667], L1[668]^L1[667] };
	assign out[331:328]   = { L1[659]^L1[662]^L1[657], L1[658]^L1[661]^L1[656]^L1[659], L1[657]^L1[660]^L1[659]^L1[663]^L1[658], L1[656]^L1[663]^L1[658] };
	assign out[327:324]   = { L1[655]^L1[650], L1[654]^L1[649], L1[653]^L1[648]^L1[651], L1[652]^L1[651] };
	assign out[323:320]   = { L1[643]^L1[646]^L1[641], L1[642]^L1[645]^L1[640]^L1[643], L1[641]^L1[644]^L1[643]^L1[647]^L1[642], L1[640]^L1[647]^L1[642] };
	assign out[319:316]   = { L1[639]^L1[634], L1[638]^L1[633], L1[637]^L1[632]^L1[635], L1[636]^L1[635] };
	assign out[315:312]   = { L1[627]^L1[630]^L1[625], L1[626]^L1[629]^L1[624]^L1[627], L1[625]^L1[628]^L1[627]^L1[631]^L1[626], L1[624]^L1[631]^L1[626] };
	assign out[311:308]   = { L1[623]^L1[618], L1[622]^L1[617], L1[621]^L1[616]^L1[619], L1[620]^L1[619] };
	assign out[307:304]   = { L1[611]^L1[614]^L1[609], L1[610]^L1[613]^L1[608]^L1[611], L1[609]^L1[612]^L1[611]^L1[615]^L1[610], L1[608]^L1[615]^L1[610] };
	assign out[303:300]   = { L1[607]^L1[602], L1[606]^L1[601], L1[605]^L1[600]^L1[603], L1[604]^L1[603] };
	assign out[299:296]   = { L1[595]^L1[598]^L1[593], L1[594]^L1[597]^L1[592]^L1[595], L1[593]^L1[596]^L1[595]^L1[599]^L1[594], L1[592]^L1[599]^L1[594] };
	assign out[295:292]   = { L1[591]^L1[586], L1[590]^L1[585], L1[589]^L1[584]^L1[587], L1[588]^L1[587] };
	assign out[291:288]   = { L1[579]^L1[582]^L1[577], L1[578]^L1[581]^L1[576]^L1[579], L1[577]^L1[580]^L1[579]^L1[583]^L1[578], L1[576]^L1[583]^L1[578] };
	assign out[287:284]   = { L1[575]^L1[570], L1[574]^L1[569], L1[573]^L1[568]^L1[571], L1[572]^L1[571] };
	assign out[283:280]   = { L1[563]^L1[566]^L1[561], L1[562]^L1[565]^L1[560]^L1[563], L1[561]^L1[564]^L1[563]^L1[567]^L1[562], L1[560]^L1[567]^L1[562] };
	assign out[279:276]   = { L1[559]^L1[554], L1[558]^L1[553], L1[557]^L1[552]^L1[555], L1[556]^L1[555] };
	assign out[275:272]   = { L1[547]^L1[550]^L1[545], L1[546]^L1[549]^L1[544]^L1[547], L1[545]^L1[548]^L1[547]^L1[551]^L1[546], L1[544]^L1[551]^L1[546] };
	assign out[271:268]   = { L1[543]^L1[538], L1[542]^L1[537], L1[541]^L1[536]^L1[539], L1[540]^L1[539] };
	assign out[267:264]   = { L1[531]^L1[534]^L1[529], L1[530]^L1[533]^L1[528]^L1[531], L1[529]^L1[532]^L1[531]^L1[535]^L1[530], L1[528]^L1[535]^L1[530] };
	assign out[263:260]   = { L1[527]^L1[522], L1[526]^L1[521], L1[525]^L1[520]^L1[523], L1[524]^L1[523] };
	assign out[259:256]   = { L1[515]^L1[518]^L1[513], L1[514]^L1[517]^L1[512]^L1[515], L1[513]^L1[516]^L1[515]^L1[519]^L1[514], L1[512]^L1[519]^L1[514] };
	assign out[255:252]   = { L1[511]^L1[506], L1[510]^L1[505], L1[509]^L1[504]^L1[507], L1[508]^L1[507] };
	assign out[251:248]   = { L1[499]^L1[502]^L1[497], L1[498]^L1[501]^L1[496]^L1[499], L1[497]^L1[500]^L1[499]^L1[503]^L1[498], L1[496]^L1[503]^L1[498] };
	assign out[247:244]   = { L1[495]^L1[490], L1[494]^L1[489], L1[493]^L1[488]^L1[491], L1[492]^L1[491] };
	assign out[243:240]   = { L1[483]^L1[486]^L1[481], L1[482]^L1[485]^L1[480]^L1[483], L1[481]^L1[484]^L1[483]^L1[487]^L1[482], L1[480]^L1[487]^L1[482] };
	assign out[239:236]   = { L1[479]^L1[474], L1[478]^L1[473], L1[477]^L1[472]^L1[475], L1[476]^L1[475] };
	assign out[235:232]   = { L1[467]^L1[470]^L1[465], L1[466]^L1[469]^L1[464]^L1[467], L1[465]^L1[468]^L1[467]^L1[471]^L1[466], L1[464]^L1[471]^L1[466] };
	assign out[231:228]   = { L1[463]^L1[458], L1[462]^L1[457], L1[461]^L1[456]^L1[459], L1[460]^L1[459] };
	assign out[227:224]   = { L1[451]^L1[454]^L1[449], L1[450]^L1[453]^L1[448]^L1[451], L1[449]^L1[452]^L1[451]^L1[455]^L1[450], L1[448]^L1[455]^L1[450] };
	assign out[223:220]   = { L1[447]^L1[442], L1[446]^L1[441], L1[445]^L1[440]^L1[443], L1[444]^L1[443] };
	assign out[219:216]   = { L1[435]^L1[438]^L1[433], L1[434]^L1[437]^L1[432]^L1[435], L1[433]^L1[436]^L1[435]^L1[439]^L1[434], L1[432]^L1[439]^L1[434] };
	assign out[215:212]   = { L1[431]^L1[426], L1[430]^L1[425], L1[429]^L1[424]^L1[427], L1[428]^L1[427] };
	assign out[211:208]   = { L1[419]^L1[422]^L1[417], L1[418]^L1[421]^L1[416]^L1[419], L1[417]^L1[420]^L1[419]^L1[423]^L1[418], L1[416]^L1[423]^L1[418] };
	assign out[207:204]   = { L1[415]^L1[410], L1[414]^L1[409], L1[413]^L1[408]^L1[411], L1[412]^L1[411] };
	assign out[203:200]   = { L1[403]^L1[406]^L1[401], L1[402]^L1[405]^L1[400]^L1[403], L1[401]^L1[404]^L1[403]^L1[407]^L1[402], L1[400]^L1[407]^L1[402] };
	assign out[199:196]   = { L1[399]^L1[394], L1[398]^L1[393], L1[397]^L1[392]^L1[395], L1[396]^L1[395] };
	assign out[195:192]   = { L1[387]^L1[390]^L1[385], L1[386]^L1[389]^L1[384]^L1[387], L1[385]^L1[388]^L1[387]^L1[391]^L1[386], L1[384]^L1[391]^L1[386] };
	assign out[191:188]   = { L1[383]^L1[378], L1[382]^L1[377], L1[381]^L1[376]^L1[379], L1[380]^L1[379] };
	assign out[187:184]   = { L1[371]^L1[374]^L1[369], L1[370]^L1[373]^L1[368]^L1[371], L1[369]^L1[372]^L1[371]^L1[375]^L1[370], L1[368]^L1[375]^L1[370] };
	assign out[183:180]   = { L1[367]^L1[362], L1[366]^L1[361], L1[365]^L1[360]^L1[363], L1[364]^L1[363] };
	assign out[179:176]   = { L1[355]^L1[358]^L1[353], L1[354]^L1[357]^L1[352]^L1[355], L1[353]^L1[356]^L1[355]^L1[359]^L1[354], L1[352]^L1[359]^L1[354] };
	assign out[175:172]   = { L1[351]^L1[346], L1[350]^L1[345], L1[349]^L1[344]^L1[347], L1[348]^L1[347] };
	assign out[171:168]   = { L1[339]^L1[342]^L1[337], L1[338]^L1[341]^L1[336]^L1[339], L1[337]^L1[340]^L1[339]^L1[343]^L1[338], L1[336]^L1[343]^L1[338] };
	assign out[167:164]   = { L1[335]^L1[330], L1[334]^L1[329], L1[333]^L1[328]^L1[331], L1[332]^L1[331] };
	assign out[163:160]   = { L1[323]^L1[326]^L1[321], L1[322]^L1[325]^L1[320]^L1[323], L1[321]^L1[324]^L1[323]^L1[327]^L1[322], L1[320]^L1[327]^L1[322] };
	assign out[159:156]   = { L1[319]^L1[314], L1[318]^L1[313], L1[317]^L1[312]^L1[315], L1[316]^L1[315] };
	assign out[155:152]   = { L1[307]^L1[310]^L1[305], L1[306]^L1[309]^L1[304]^L1[307], L1[305]^L1[308]^L1[307]^L1[311]^L1[306], L1[304]^L1[311]^L1[306] };
	assign out[151:148]   = { L1[303]^L1[298], L1[302]^L1[297], L1[301]^L1[296]^L1[299], L1[300]^L1[299] };
	assign out[147:144]   = { L1[291]^L1[294]^L1[289], L1[290]^L1[293]^L1[288]^L1[291], L1[289]^L1[292]^L1[291]^L1[295]^L1[290], L1[288]^L1[295]^L1[290] };
	assign out[143:140]   = { L1[287]^L1[282], L1[286]^L1[281], L1[285]^L1[280]^L1[283], L1[284]^L1[283] };
	assign out[139:136]   = { L1[275]^L1[278]^L1[273], L1[274]^L1[277]^L1[272]^L1[275], L1[273]^L1[276]^L1[275]^L1[279]^L1[274], L1[272]^L1[279]^L1[274] };
	assign out[135:132]   = { L1[271]^L1[266], L1[270]^L1[265], L1[269]^L1[264]^L1[267], L1[268]^L1[267] };
	assign out[131:128]   = { L1[259]^L1[262]^L1[257], L1[258]^L1[261]^L1[256]^L1[259], L1[257]^L1[260]^L1[259]^L1[263]^L1[258], L1[256]^L1[263]^L1[258] };
	assign out[127:124]   = { L1[255]^L1[250], L1[254]^L1[249], L1[253]^L1[248]^L1[251], L1[252]^L1[251] };
	assign out[123:120]   = { L1[243]^L1[246]^L1[241], L1[242]^L1[245]^L1[240]^L1[243], L1[241]^L1[244]^L1[243]^L1[247]^L1[242], L1[240]^L1[247]^L1[242] };
	assign out[119:116]   = { L1[239]^L1[234], L1[238]^L1[233], L1[237]^L1[232]^L1[235], L1[236]^L1[235] };
	assign out[115:112]   = { L1[227]^L1[230]^L1[225], L1[226]^L1[229]^L1[224]^L1[227], L1[225]^L1[228]^L1[227]^L1[231]^L1[226], L1[224]^L1[231]^L1[226] };
	assign out[111:108]   = { L1[223]^L1[218], L1[222]^L1[217], L1[221]^L1[216]^L1[219], L1[220]^L1[219] };
	assign out[107:104]   = { L1[211]^L1[214]^L1[209], L1[210]^L1[213]^L1[208]^L1[211], L1[209]^L1[212]^L1[211]^L1[215]^L1[210], L1[208]^L1[215]^L1[210] };
	assign out[103:100]   = { L1[207]^L1[202], L1[206]^L1[201], L1[205]^L1[200]^L1[203], L1[204]^L1[203] };
	assign out[ 99: 96]   = { L1[195]^L1[198]^L1[193], L1[194]^L1[197]^L1[192]^L1[195], L1[193]^L1[196]^L1[195]^L1[199]^L1[194], L1[192]^L1[199]^L1[194] };
	assign out[ 95: 92]   = { L1[191]^L1[186], L1[190]^L1[185], L1[189]^L1[184]^L1[187], L1[188]^L1[187] };
	assign out[ 91: 88]   = { L1[179]^L1[182]^L1[177], L1[178]^L1[181]^L1[176]^L1[179], L1[177]^L1[180]^L1[179]^L1[183]^L1[178], L1[176]^L1[183]^L1[178] };
	assign out[ 87: 84]   = { L1[175]^L1[170], L1[174]^L1[169], L1[173]^L1[168]^L1[171], L1[172]^L1[171] };
	assign out[ 83: 80]   = { L1[163]^L1[166]^L1[161], L1[162]^L1[165]^L1[160]^L1[163], L1[161]^L1[164]^L1[163]^L1[167]^L1[162], L1[160]^L1[167]^L1[162] };
	assign out[ 79: 76]   = { L1[159]^L1[154], L1[158]^L1[153], L1[157]^L1[152]^L1[155], L1[156]^L1[155] };
	assign out[ 75: 72]   = { L1[147]^L1[150]^L1[145], L1[146]^L1[149]^L1[144]^L1[147], L1[145]^L1[148]^L1[147]^L1[151]^L1[146], L1[144]^L1[151]^L1[146] };
	assign out[ 71: 68]   = { L1[143]^L1[138], L1[142]^L1[137], L1[141]^L1[136]^L1[139], L1[140]^L1[139] };
	assign out[ 67: 64]   = { L1[131]^L1[134]^L1[129], L1[130]^L1[133]^L1[128]^L1[131], L1[129]^L1[132]^L1[131]^L1[135]^L1[130], L1[128]^L1[135]^L1[130] };
	assign out[ 63: 60]   = { L1[127]^L1[122], L1[126]^L1[121], L1[125]^L1[120]^L1[123], L1[124]^L1[123] };
	assign out[ 59: 56]   = { L1[115]^L1[118]^L1[113], L1[114]^L1[117]^L1[112]^L1[115], L1[113]^L1[116]^L1[115]^L1[119]^L1[114], L1[112]^L1[119]^L1[114] };
	assign out[ 55: 52]   = { L1[111]^L1[106], L1[110]^L1[105], L1[109]^L1[104]^L1[107], L1[108]^L1[107] };
	assign out[ 51: 48]   = { L1[99]^L1[102]^L1[97], L1[98]^L1[101]^L1[96]^L1[99], L1[97]^L1[100]^L1[99]^L1[103]^L1[98], L1[96]^L1[103]^L1[98] };
	assign out[ 47: 44]   = { L1[95]^L1[90], L1[94]^L1[89], L1[93]^L1[88]^L1[91], L1[92]^L1[91] };
	assign out[ 43: 40]   = { L1[83]^L1[86]^L1[81], L1[82]^L1[85]^L1[80]^L1[83], L1[81]^L1[84]^L1[83]^L1[87]^L1[82], L1[80]^L1[87]^L1[82] };
	assign out[ 39: 36]   = { L1[79]^L1[74], L1[78]^L1[73], L1[77]^L1[72]^L1[75], L1[76]^L1[75] };
	assign out[ 35: 32]   = { L1[67]^L1[70]^L1[65], L1[66]^L1[69]^L1[64]^L1[67], L1[65]^L1[68]^L1[67]^L1[71]^L1[66], L1[64]^L1[71]^L1[66] };
	assign out[ 31: 28]   = { L1[63]^L1[58], L1[62]^L1[57], L1[61]^L1[56]^L1[59], L1[60]^L1[59] };
	assign out[ 27: 24]   = { L1[51]^L1[54]^L1[49], L1[50]^L1[53]^L1[48]^L1[51], L1[49]^L1[52]^L1[51]^L1[55]^L1[50], L1[48]^L1[55]^L1[50] };
	assign out[ 23: 20]   = { L1[47]^L1[42], L1[46]^L1[41], L1[45]^L1[40]^L1[43], L1[44]^L1[43] };
	assign out[ 19: 16]   = { L1[35]^L1[38]^L1[33], L1[34]^L1[37]^L1[32]^L1[35], L1[33]^L1[36]^L1[35]^L1[39]^L1[34], L1[32]^L1[39]^L1[34] };
	assign out[ 15: 12]   = { L1[31]^L1[26], L1[30]^L1[25], L1[29]^L1[24]^L1[27], L1[28]^L1[27] };
	assign out[ 11:  8]   = { L1[19]^L1[22]^L1[17], L1[18]^L1[21]^L1[16]^L1[19], L1[17]^L1[20]^L1[19]^L1[23]^L1[18], L1[16]^L1[23]^L1[18] };
	assign out[  7:  4]   = { L1[15]^L1[10], L1[14]^L1[9], L1[13]^L1[8]^L1[11], L1[12]^L1[11] };
	assign out[  3:  0]   = { L1[3]^L1[6]^L1[1], L1[2]^L1[5]^L1[0]^L1[3], L1[1]^L1[4]^L1[3]^L1[7]^L1[2], L1[0]^L1[7]^L1[2] };

endmodule 

