module jh_final (
	input [1023:0] in,
	output [1023:0] out
);

	 assign { out[7], out[263], out[519], out[775] } = in[3:0];
	 assign { out[6], out[262], out[518], out[774] } = in[11:8];
	 assign { out[5], out[261], out[517], out[773] } = in[19:16];
	 assign { out[4], out[260], out[516], out[772] } = in[27:24];
	 assign { out[3], out[259], out[515], out[771] } = in[35:32];
	 assign { out[2], out[258], out[514], out[770] } = in[43:40];
	 assign { out[1], out[257], out[513], out[769] } = in[51:48];
	 assign { out[0], out[256], out[512], out[768] } = in[59:56];
	 assign { out[15], out[271], out[527], out[783] } = in[67:64];
	 assign { out[14], out[270], out[526], out[782] } = in[75:72];
	 assign { out[13], out[269], out[525], out[781] } = in[83:80];
	 assign { out[12], out[268], out[524], out[780] } = in[91:88];
	 assign { out[11], out[267], out[523], out[779] } = in[99:96];
	 assign { out[10], out[266], out[522], out[778] } = in[107:104];
	 assign { out[9], out[265], out[521], out[777] } = in[115:112];
	 assign { out[8], out[264], out[520], out[776] } = in[123:120];
	 assign { out[23], out[279], out[535], out[791] } = in[131:128];
	 assign { out[22], out[278], out[534], out[790] } = in[139:136];
	 assign { out[21], out[277], out[533], out[789] } = in[147:144];
	 assign { out[20], out[276], out[532], out[788] } = in[155:152];
	 assign { out[19], out[275], out[531], out[787] } = in[163:160];
	 assign { out[18], out[274], out[530], out[786] } = in[171:168];
	 assign { out[17], out[273], out[529], out[785] } = in[179:176];
	 assign { out[16], out[272], out[528], out[784] } = in[187:184];
	 assign { out[31], out[287], out[543], out[799] } = in[195:192];
	 assign { out[30], out[286], out[542], out[798] } = in[203:200];
	 assign { out[29], out[285], out[541], out[797] } = in[211:208];
	 assign { out[28], out[284], out[540], out[796] } = in[219:216];
	 assign { out[27], out[283], out[539], out[795] } = in[227:224];
	 assign { out[26], out[282], out[538], out[794] } = in[235:232];
	 assign { out[25], out[281], out[537], out[793] } = in[243:240];
	 assign { out[24], out[280], out[536], out[792] } = in[251:248];
	 assign { out[39], out[295], out[551], out[807] } = in[259:256];
	 assign { out[38], out[294], out[550], out[806] } = in[267:264];
	 assign { out[37], out[293], out[549], out[805] } = in[275:272];
	 assign { out[36], out[292], out[548], out[804] } = in[283:280];
	 assign { out[35], out[291], out[547], out[803] } = in[291:288];
	 assign { out[34], out[290], out[546], out[802] } = in[299:296];
	 assign { out[33], out[289], out[545], out[801] } = in[307:304];
	 assign { out[32], out[288], out[544], out[800] } = in[315:312];
	 assign { out[47], out[303], out[559], out[815] } = in[323:320];
	 assign { out[46], out[302], out[558], out[814] } = in[331:328];
	 assign { out[45], out[301], out[557], out[813] } = in[339:336];
	 assign { out[44], out[300], out[556], out[812] } = in[347:344];
	 assign { out[43], out[299], out[555], out[811] } = in[355:352];
	 assign { out[42], out[298], out[554], out[810] } = in[363:360];
	 assign { out[41], out[297], out[553], out[809] } = in[371:368];
	 assign { out[40], out[296], out[552], out[808] } = in[379:376];
	 assign { out[55], out[311], out[567], out[823] } = in[387:384];
	 assign { out[54], out[310], out[566], out[822] } = in[395:392];
	 assign { out[53], out[309], out[565], out[821] } = in[403:400];
	 assign { out[52], out[308], out[564], out[820] } = in[411:408];
	 assign { out[51], out[307], out[563], out[819] } = in[419:416];
	 assign { out[50], out[306], out[562], out[818] } = in[427:424];
	 assign { out[49], out[305], out[561], out[817] } = in[435:432];
	 assign { out[48], out[304], out[560], out[816] } = in[443:440];
	 assign { out[63], out[319], out[575], out[831] } = in[451:448];
	 assign { out[62], out[318], out[574], out[830] } = in[459:456];
	 assign { out[61], out[317], out[573], out[829] } = in[467:464];
	 assign { out[60], out[316], out[572], out[828] } = in[475:472];
	 assign { out[59], out[315], out[571], out[827] } = in[483:480];
	 assign { out[58], out[314], out[570], out[826] } = in[491:488];
	 assign { out[57], out[313], out[569], out[825] } = in[499:496];
	 assign { out[56], out[312], out[568], out[824] } = in[507:504];
	 assign { out[71], out[327], out[583], out[839] } = in[515:512];
	 assign { out[70], out[326], out[582], out[838] } = in[523:520];
	 assign { out[69], out[325], out[581], out[837] } = in[531:528];
	 assign { out[68], out[324], out[580], out[836] } = in[539:536];
	 assign { out[67], out[323], out[579], out[835] } = in[547:544];
	 assign { out[66], out[322], out[578], out[834] } = in[555:552];
	 assign { out[65], out[321], out[577], out[833] } = in[563:560];
	 assign { out[64], out[320], out[576], out[832] } = in[571:568];
	 assign { out[79], out[335], out[591], out[847] } = in[579:576];
	 assign { out[78], out[334], out[590], out[846] } = in[587:584];
	 assign { out[77], out[333], out[589], out[845] } = in[595:592];
	 assign { out[76], out[332], out[588], out[844] } = in[603:600];
	 assign { out[75], out[331], out[587], out[843] } = in[611:608];
	 assign { out[74], out[330], out[586], out[842] } = in[619:616];
	 assign { out[73], out[329], out[585], out[841] } = in[627:624];
	 assign { out[72], out[328], out[584], out[840] } = in[635:632];
	 assign { out[87], out[343], out[599], out[855] } = in[643:640];
	 assign { out[86], out[342], out[598], out[854] } = in[651:648];
	 assign { out[85], out[341], out[597], out[853] } = in[659:656];
	 assign { out[84], out[340], out[596], out[852] } = in[667:664];
	 assign { out[83], out[339], out[595], out[851] } = in[675:672];
	 assign { out[82], out[338], out[594], out[850] } = in[683:680];
	 assign { out[81], out[337], out[593], out[849] } = in[691:688];
	 assign { out[80], out[336], out[592], out[848] } = in[699:696];
	 assign { out[95], out[351], out[607], out[863] } = in[707:704];
	 assign { out[94], out[350], out[606], out[862] } = in[715:712];
	 assign { out[93], out[349], out[605], out[861] } = in[723:720];
	 assign { out[92], out[348], out[604], out[860] } = in[731:728];
	 assign { out[91], out[347], out[603], out[859] } = in[739:736];
	 assign { out[90], out[346], out[602], out[858] } = in[747:744];
	 assign { out[89], out[345], out[601], out[857] } = in[755:752];
	 assign { out[88], out[344], out[600], out[856] } = in[763:760];
	 assign { out[103], out[359], out[615], out[871] } = in[771:768];
	 assign { out[102], out[358], out[614], out[870] } = in[779:776];
	 assign { out[101], out[357], out[613], out[869] } = in[787:784];
	 assign { out[100], out[356], out[612], out[868] } = in[795:792];
	 assign { out[99], out[355], out[611], out[867] } = in[803:800];
	 assign { out[98], out[354], out[610], out[866] } = in[811:808];
	 assign { out[97], out[353], out[609], out[865] } = in[819:816];
	 assign { out[96], out[352], out[608], out[864] } = in[827:824];
	 assign { out[111], out[367], out[623], out[879] } = in[835:832];
	 assign { out[110], out[366], out[622], out[878] } = in[843:840];
	 assign { out[109], out[365], out[621], out[877] } = in[851:848];
	 assign { out[108], out[364], out[620], out[876] } = in[859:856];
	 assign { out[107], out[363], out[619], out[875] } = in[867:864];
	 assign { out[106], out[362], out[618], out[874] } = in[875:872];
	 assign { out[105], out[361], out[617], out[873] } = in[883:880];
	 assign { out[104], out[360], out[616], out[872] } = in[891:888];
	 assign { out[119], out[375], out[631], out[887] } = in[899:896];
	 assign { out[118], out[374], out[630], out[886] } = in[907:904];
	 assign { out[117], out[373], out[629], out[885] } = in[915:912];
	 assign { out[116], out[372], out[628], out[884] } = in[923:920];
	 assign { out[115], out[371], out[627], out[883] } = in[931:928];
	 assign { out[114], out[370], out[626], out[882] } = in[939:936];
	 assign { out[113], out[369], out[625], out[881] } = in[947:944];
	 assign { out[112], out[368], out[624], out[880] } = in[955:952];
	 assign { out[127], out[383], out[639], out[895] } = in[963:960];
	 assign { out[126], out[382], out[638], out[894] } = in[971:968];
	 assign { out[125], out[381], out[637], out[893] } = in[979:976];
	 assign { out[124], out[380], out[636], out[892] } = in[987:984];
	 assign { out[123], out[379], out[635], out[891] } = in[995:992];
	 assign { out[122], out[378], out[634], out[890] } = in[1003:1000];
	 assign { out[121], out[377], out[633], out[889] } = in[1011:1008];
	 assign { out[120], out[376], out[632], out[888] } = in[1019:1016];
	 assign { out[135], out[391], out[647], out[903] } = in[7:4];
	 assign { out[134], out[390], out[646], out[902] } = in[15:12];
	 assign { out[133], out[389], out[645], out[901] } = in[23:20];
	 assign { out[132], out[388], out[644], out[900] } = in[31:28];
	 assign { out[131], out[387], out[643], out[899] } = in[39:36];
	 assign { out[130], out[386], out[642], out[898] } = in[47:44];
	 assign { out[129], out[385], out[641], out[897] } = in[55:52];
	 assign { out[128], out[384], out[640], out[896] } = in[63:60];
	 assign { out[143], out[399], out[655], out[911] } = in[71:68];
	 assign { out[142], out[398], out[654], out[910] } = in[79:76];
	 assign { out[141], out[397], out[653], out[909] } = in[87:84];
	 assign { out[140], out[396], out[652], out[908] } = in[95:92];
	 assign { out[139], out[395], out[651], out[907] } = in[103:100];
	 assign { out[138], out[394], out[650], out[906] } = in[111:108];
	 assign { out[137], out[393], out[649], out[905] } = in[119:116];
	 assign { out[136], out[392], out[648], out[904] } = in[127:124];
	 assign { out[151], out[407], out[663], out[919] } = in[135:132];
	 assign { out[150], out[406], out[662], out[918] } = in[143:140];
	 assign { out[149], out[405], out[661], out[917] } = in[151:148];
	 assign { out[148], out[404], out[660], out[916] } = in[159:156];
	 assign { out[147], out[403], out[659], out[915] } = in[167:164];
	 assign { out[146], out[402], out[658], out[914] } = in[175:172];
	 assign { out[145], out[401], out[657], out[913] } = in[183:180];
	 assign { out[144], out[400], out[656], out[912] } = in[191:188];
	 assign { out[159], out[415], out[671], out[927] } = in[199:196];
	 assign { out[158], out[414], out[670], out[926] } = in[207:204];
	 assign { out[157], out[413], out[669], out[925] } = in[215:212];
	 assign { out[156], out[412], out[668], out[924] } = in[223:220];
	 assign { out[155], out[411], out[667], out[923] } = in[231:228];
	 assign { out[154], out[410], out[666], out[922] } = in[239:236];
	 assign { out[153], out[409], out[665], out[921] } = in[247:244];
	 assign { out[152], out[408], out[664], out[920] } = in[255:252];
	 assign { out[167], out[423], out[679], out[935] } = in[263:260];
	 assign { out[166], out[422], out[678], out[934] } = in[271:268];
	 assign { out[165], out[421], out[677], out[933] } = in[279:276];
	 assign { out[164], out[420], out[676], out[932] } = in[287:284];
	 assign { out[163], out[419], out[675], out[931] } = in[295:292];
	 assign { out[162], out[418], out[674], out[930] } = in[303:300];
	 assign { out[161], out[417], out[673], out[929] } = in[311:308];
	 assign { out[160], out[416], out[672], out[928] } = in[319:316];
	 assign { out[175], out[431], out[687], out[943] } = in[327:324];
	 assign { out[174], out[430], out[686], out[942] } = in[335:332];
	 assign { out[173], out[429], out[685], out[941] } = in[343:340];
	 assign { out[172], out[428], out[684], out[940] } = in[351:348];
	 assign { out[171], out[427], out[683], out[939] } = in[359:356];
	 assign { out[170], out[426], out[682], out[938] } = in[367:364];
	 assign { out[169], out[425], out[681], out[937] } = in[375:372];
	 assign { out[168], out[424], out[680], out[936] } = in[383:380];
	 assign { out[183], out[439], out[695], out[951] } = in[391:388];
	 assign { out[182], out[438], out[694], out[950] } = in[399:396];
	 assign { out[181], out[437], out[693], out[949] } = in[407:404];
	 assign { out[180], out[436], out[692], out[948] } = in[415:412];
	 assign { out[179], out[435], out[691], out[947] } = in[423:420];
	 assign { out[178], out[434], out[690], out[946] } = in[431:428];
	 assign { out[177], out[433], out[689], out[945] } = in[439:436];
	 assign { out[176], out[432], out[688], out[944] } = in[447:444];
	 assign { out[191], out[447], out[703], out[959] } = in[455:452];
	 assign { out[190], out[446], out[702], out[958] } = in[463:460];
	 assign { out[189], out[445], out[701], out[957] } = in[471:468];
	 assign { out[188], out[444], out[700], out[956] } = in[479:476];
	 assign { out[187], out[443], out[699], out[955] } = in[487:484];
	 assign { out[186], out[442], out[698], out[954] } = in[495:492];
	 assign { out[185], out[441], out[697], out[953] } = in[503:500];
	 assign { out[184], out[440], out[696], out[952] } = in[511:508];
	 assign { out[199], out[455], out[711], out[967] } = in[519:516];
	 assign { out[198], out[454], out[710], out[966] } = in[527:524];
	 assign { out[197], out[453], out[709], out[965] } = in[535:532];
	 assign { out[196], out[452], out[708], out[964] } = in[543:540];
	 assign { out[195], out[451], out[707], out[963] } = in[551:548];
	 assign { out[194], out[450], out[706], out[962] } = in[559:556];
	 assign { out[193], out[449], out[705], out[961] } = in[567:564];
	 assign { out[192], out[448], out[704], out[960] } = in[575:572];
	 assign { out[207], out[463], out[719], out[975] } = in[583:580];
	 assign { out[206], out[462], out[718], out[974] } = in[591:588];
	 assign { out[205], out[461], out[717], out[973] } = in[599:596];
	 assign { out[204], out[460], out[716], out[972] } = in[607:604];
	 assign { out[203], out[459], out[715], out[971] } = in[615:612];
	 assign { out[202], out[458], out[714], out[970] } = in[623:620];
	 assign { out[201], out[457], out[713], out[969] } = in[631:628];
	 assign { out[200], out[456], out[712], out[968] } = in[639:636];
	 assign { out[215], out[471], out[727], out[983] } = in[647:644];
	 assign { out[214], out[470], out[726], out[982] } = in[655:652];
	 assign { out[213], out[469], out[725], out[981] } = in[663:660];
	 assign { out[212], out[468], out[724], out[980] } = in[671:668];
	 assign { out[211], out[467], out[723], out[979] } = in[679:676];
	 assign { out[210], out[466], out[722], out[978] } = in[687:684];
	 assign { out[209], out[465], out[721], out[977] } = in[695:692];
	 assign { out[208], out[464], out[720], out[976] } = in[703:700];
	 assign { out[223], out[479], out[735], out[991] } = in[711:708];
	 assign { out[222], out[478], out[734], out[990] } = in[719:716];
	 assign { out[221], out[477], out[733], out[989] } = in[727:724];
	 assign { out[220], out[476], out[732], out[988] } = in[735:732];
	 assign { out[219], out[475], out[731], out[987] } = in[743:740];
	 assign { out[218], out[474], out[730], out[986] } = in[751:748];
	 assign { out[217], out[473], out[729], out[985] } = in[759:756];
	 assign { out[216], out[472], out[728], out[984] } = in[767:764];
	 assign { out[231], out[487], out[743], out[999] } = in[775:772];
	 assign { out[230], out[486], out[742], out[998] } = in[783:780];
	 assign { out[229], out[485], out[741], out[997] } = in[791:788];
	 assign { out[228], out[484], out[740], out[996] } = in[799:796];
	 assign { out[227], out[483], out[739], out[995] } = in[807:804];
	 assign { out[226], out[482], out[738], out[994] } = in[815:812];
	 assign { out[225], out[481], out[737], out[993] } = in[823:820];
	 assign { out[224], out[480], out[736], out[992] } = in[831:828];
	 assign { out[239], out[495], out[751], out[1007] } = in[839:836];
	 assign { out[238], out[494], out[750], out[1006] } = in[847:844];
	 assign { out[237], out[493], out[749], out[1005] } = in[855:852];
	 assign { out[236], out[492], out[748], out[1004] } = in[863:860];
	 assign { out[235], out[491], out[747], out[1003] } = in[871:868];
	 assign { out[234], out[490], out[746], out[1002] } = in[879:876];
	 assign { out[233], out[489], out[745], out[1001] } = in[887:884];
	 assign { out[232], out[488], out[744], out[1000] } = in[895:892];
	 assign { out[247], out[503], out[759], out[1015] } = in[903:900];
	 assign { out[246], out[502], out[758], out[1014] } = in[911:908];
	 assign { out[245], out[501], out[757], out[1013] } = in[919:916];
	 assign { out[244], out[500], out[756], out[1012] } = in[927:924];
	 assign { out[243], out[499], out[755], out[1011] } = in[935:932];
	 assign { out[242], out[498], out[754], out[1010] } = in[943:940];
	 assign { out[241], out[497], out[753], out[1009] } = in[951:948];
	 assign { out[240], out[496], out[752], out[1008] } = in[959:956];
	 assign { out[255], out[511], out[767], out[1023] } = in[967:964];
	 assign { out[254], out[510], out[766], out[1022] } = in[975:972];
	 assign { out[253], out[509], out[765], out[1021] } = in[983:980];
	 assign { out[252], out[508], out[764], out[1020] } = in[991:988];
	 assign { out[251], out[507], out[763], out[1019] } = in[999:996];
	 assign { out[250], out[506], out[762], out[1018] } = in[1007:1004];
	 assign { out[249], out[505], out[761], out[1017] } = in[1015:1012];
	 assign { out[248], out[504], out[760], out[1016] } = in[1023:1020];

endmodule

